`timescale 1ns / 1ps
`include "all_cmos_tf_rst_mnist.v"
`include "all_cmos_tf_rst.v"

module mnist_neural_network(
    input wire clk,
    input wire rst,
    input wire [115:0] input_layer, // TODO: widen if needed
    output wire [255:0] Z
);

  // Internal signals
  wire [255:0] Y; // layer 1 outputs feed layer 3

  // instantiate function_0 for neuron0_1
  function_0 neuron0_1 (
      .a(~input_layer[871]),
      .b(~input_layer[385]),
      .c(~input_layer[330]),
      .d(~input_layer[918]),
      .e(~input_layer[1216]),
      .y(Y[0]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1_1
  function_1 neuron1_1 (
      .a(~input_layer[302]),
      .b(~input_layer[367]),
      .c(~input_layer[320]),
      .d(input_layer[460]),
      .y(Y[1]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_2 for neuron2_1
  function_2 neuron2_1 (
      .a(input_layer[1200]),
      .b(input_layer[837]),
      .c(~input_layer[1413]),
      .d(input_layer[670]),
      .e(input_layer[103]),
      .f(input_layer[1556]),
      .y(Y[2]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron3_1
  function_3 neuron3_1 (
      .a(~input_layer[417]),
      .b(~input_layer[1241]),
      .c(~input_layer[1058]),
      .d(~input_layer[600]),
      .y(Y[3]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron4_1
  function_4 neuron4_1 (
      .a(~input_layer[913]),
      .b(~input_layer[301]),
      .c(~input_layer[1242]),
      .d(~input_layer[1382]),
      .e(~input_layer[116]),
      .y(Y[4]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron5_1
  function_5 neuron5_1 (
      .a(~input_layer[330]),
      .b(~input_layer[969]),
      .c(input_layer[815]),
      .d(~input_layer[465]),
      .e(~input_layer[375]),
      .f(input_layer[233]),
      .y(Y[5]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron6_1
  function_6 neuron6_1 (
      .a(~input_layer[587]),
      .b(~input_layer[1210]),
      .c(input_layer[1228]),
      .d(input_layer[1242]),
      .e(input_layer[224]),
      .f(~input_layer[952]),
      .y(Y[6]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron7_1
  function_3 neuron7_1 (
      .a(~input_layer[459]),
      .b(input_layer[1027]),
      .c(~input_layer[1068]),
      .d(~input_layer[453]),
      .y(Y[7]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron8_1
  function_7 neuron8_1 (
      .a(input_layer[1020]),
      .b(~input_layer[733]),
      .c(input_layer[95]),
      .d(input_layer[1321]),
      .y(Y[8]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron9_1
  function_8 neuron9_1 (
      .a(input_layer[201]),
      .b(~input_layer[862]),
      .c(input_layer[1362]),
      .d(input_layer[459]),
      .y(Y[9]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_9 for neuron10_1
  function_9 neuron10_1 (
      .a(input_layer[968]),
      .b(input_layer[133]),
      .c(~input_layer[1268]),
      .d(input_layer[942]),
      .e(input_layer[1338]),
      .f(~input_layer[931]),
      .y(Y[10]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron11_1
  function_10 neuron11_1 (
      .a(~input_layer[801]),
      .b(input_layer[147]),
      .c(input_layer[517]),
      .d(~input_layer[1040]),
      .e(input_layer[559]),
      .f(~input_layer[12]),
      .y(Y[11]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron12_1
  function_3 neuron12_1 (
      .a(~input_layer[936]),
      .b(~input_layer[523]),
      .c(~input_layer[1311]),
      .d(~input_layer[847]),
      .y(Y[12]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron13_1
  function_11 neuron13_1 (
      .a(~input_layer[1275]),
      .b(input_layer[1413]),
      .c(~input_layer[428]),
      .d(~input_layer[235]),
      .y(Y[13]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron14_1
  function_12 neuron14_1 (
      .a(input_layer[773]),
      .b(~input_layer[638]),
      .c(~input_layer[746]),
      .y(Y[14]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron15_1
  function_11 neuron15_1 (
      .a(~input_layer[926]),
      .b(~input_layer[645]),
      .c(input_layer[656]),
      .d(~input_layer[303]),
      .y(Y[15]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron16_1
  function_13 neuron16_1 (
      .a(~input_layer[697]),
      .b(input_layer[791]),
      .c(~input_layer[855]),
      .d(~input_layer[333]),
      .y(Y[16]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron17_1
  function_14 neuron17_1 (
      .a(~input_layer[867]),
      .b(input_layer[1004]),
      .c(input_layer[1524]),
      .d(input_layer[1349]),
      .e(~input_layer[435]),
      .f(~input_layer[632]),
      .y(Y[17]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_15 for neuron18_1
  function_15 neuron18_1 (
      .a(input_layer[440]),
      .b(input_layer[383]),
      .c(~input_layer[480]),
      .d(~input_layer[1487]),
      .e(~input_layer[760]),
      .f(~input_layer[105]),
      .y(Y[18]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron19_1
  function_16 neuron19_1 (
      .a(input_layer[611]),
      .b(~input_layer[1084]),
      .y(Y[19]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron20_1
  function_17 neuron20_1 (
      .a(input_layer[1189]),
      .b(input_layer[445]),
      .c(~input_layer[1208]),
      .y(Y[20]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron21_1
  function_18 neuron21_1 (
      .a(input_layer[945]),
      .b(~input_layer[604]),
      .c(~input_layer[1269]),
      .d(~input_layer[1393]),
      .e(input_layer[1037]),
      .y(Y[21]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron22_1
  function_3 neuron22_1 (
      .a(~input_layer[1333]),
      .b(~input_layer[438]),
      .c(input_layer[516]),
      .d(~input_layer[143]),
      .y(Y[22]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron23_1
  function_19 neuron23_1 (
      .a(~input_layer[1442]),
      .b(~input_layer[1130]),
      .c(~input_layer[1248]),
      .d(input_layer[215]),
      .y(Y[23]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron24_1
  function_20 neuron24_1 (
      .a(~input_layer[439]),
      .b(~input_layer[852]),
      .c(input_layer[781]),
      .d(input_layer[536]),
      .e(~input_layer[174]),
      .y(Y[24]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron25_1
  function_21 neuron25_1 (
      .a(input_layer[322]),
      .b(~input_layer[482]),
      .c(input_layer[850]),
      .d(input_layer[1204]),
      .e(~input_layer[116]),
      .y(Y[25]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_22 for neuron26_1
  function_22 neuron26_1 (
      .a(input_layer[499]),
      .b(~input_layer[528]),
      .c(input_layer[376]),
      .d(input_layer[893]),
      .e(~input_layer[1525]),
      .f(~input_layer[1380]),
      .y(Y[26]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_23 for neuron27_1
  function_23 neuron27_1 (
      .a(~input_layer[621]),
      .b(input_layer[1442]),
      .c(~input_layer[1550]),
      .d(~input_layer[1558]),
      .e(input_layer[20]),
      .f(~input_layer[37]),
      .y(Y[27]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron28_1
  function_3 neuron28_1 (
      .a(~input_layer[539]),
      .b(~input_layer[1014]),
      .c(~input_layer[437]),
      .d(input_layer[1046]),
      .y(Y[28]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron29_1
  function_24 neuron29_1 (
      .a(~input_layer[775]),
      .b(input_layer[603]),
      .c(input_layer[592]),
      .y(Y[29]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron30_1
  function_1 neuron30_1 (
      .a(~input_layer[590]),
      .b(input_layer[740]),
      .c(~input_layer[1252]),
      .d(~input_layer[506]),
      .y(Y[30]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron31_1
  function_25 neuron31_1 (
      .a(input_layer[1473]),
      .b(input_layer[135]),
      .c(~input_layer[696]),
      .d(~input_layer[808]),
      .e(~input_layer[502]),
      .y(Y[31]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron32_1
  function_26 neuron32_1 (
      .a(input_layer[1277]),
      .y(Y[32]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron33_1
  function_26 neuron33_1 (
      .a(~input_layer[435]),
      .y(Y[33]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron34_1
  function_27 neuron34_1 (
      .a(~input_layer[757]),
      .b(~input_layer[923]),
      .c(~input_layer[1015]),
      .y(Y[34]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron35_1
  function_28 neuron35_1 (
      .a(~input_layer[973]),
      .b(~input_layer[432]),
      .c(~input_layer[1189]),
      .d(~input_layer[328]),
      .e(~input_layer[1213]),
      .f(~input_layer[1422]),
      .y(Y[35]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron36_1
  function_24 neuron36_1 (
      .a(~input_layer[924]),
      .b(input_layer[762]),
      .c(~input_layer[379]),
      .y(Y[36]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron37_1
  function_29 neuron37_1 (
      .a(~input_layer[660]),
      .b(input_layer[321]),
      .y(Y[37]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron38_1
  function_30 neuron38_1 (
      .a(input_layer[1435]),
      .b(input_layer[484]),
      .c(input_layer[1297]),
      .d(~input_layer[863]),
      .y(Y[38]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_15 for neuron39_1
  function_15 neuron39_1 (
      .a(input_layer[931]),
      .b(input_layer[517]),
      .c(input_layer[799]),
      .d(input_layer[1533]),
      .e(~input_layer[421]),
      .f(input_layer[505]),
      .y(Y[39]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron40_1
  function_17 neuron40_1 (
      .a(input_layer[1160]),
      .b(input_layer[376]),
      .c(input_layer[93]),
      .y(Y[40]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[41] = 1'b1;

  // instantiate function_0 for neuron42_1
  function_0 neuron42_1 (
      .a(~input_layer[488]),
      .b(~input_layer[430]),
      .c(~input_layer[583]),
      .d(~input_layer[847]),
      .e(~input_layer[1408]),
      .y(Y[42]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron43_1
  function_31 neuron43_1 (
      .a(input_layer[867]),
      .b(~input_layer[600]),
      .c(~input_layer[509]),
      .d(~input_layer[436]),
      .y(Y[43]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron44_1
  function_32 neuron44_1 (
      .a(~input_layer[1077]),
      .b(input_layer[1549]),
      .c(~input_layer[1221]),
      .d(input_layer[349]),
      .e(input_layer[1445]),
      .f(~input_layer[1451]),
      .y(Y[44]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron45_1
  function_3 neuron45_1 (
      .a(~input_layer[1102]),
      .b(~input_layer[1165]),
      .c(~input_layer[568]),
      .d(input_layer[979]),
      .y(Y[45]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron46_1
  function_8 neuron46_1 (
      .a(input_layer[1077]),
      .b(input_layer[143]),
      .c(~input_layer[1548]),
      .d(input_layer[443]),
      .y(Y[46]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron47_1
  function_21 neuron47_1 (
      .a(~input_layer[1313]),
      .b(input_layer[1442]),
      .c(input_layer[1331]),
      .d(input_layer[250]),
      .e(~input_layer[1303]),
      .y(Y[47]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron48_1
  function_33 neuron48_1 (
      .a(~input_layer[1046]),
      .b(input_layer[563]),
      .c(input_layer[1142]),
      .d(~input_layer[415]),
      .e(~input_layer[309]),
      .f(~input_layer[108]),
      .y(Y[48]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron49_1
  function_27 neuron49_1 (
      .a(~input_layer[424]),
      .b(~input_layer[1225]),
      .c(~input_layer[1350]),
      .y(Y[49]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron50_1
  function_27 neuron50_1 (
      .a(~input_layer[252]),
      .b(~input_layer[498]),
      .c(~input_layer[1181]),
      .y(Y[50]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[51] = 1'b1;

  // instantiate function_34 for neuron52_1
  function_34 neuron52_1 (
      .a(~input_layer[910]),
      .b(input_layer[1392]),
      .c(~input_layer[545]),
      .d(~input_layer[1128]),
      .e(input_layer[692]),
      .f(~input_layer[417]),
      .y(Y[52]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron53_1
  function_35 neuron53_1 (
      .a(~input_layer[1074]),
      .b(~input_layer[1206]),
      .c(~input_layer[1263]),
      .d(input_layer[1417]),
      .e(input_layer[452]),
      .y(Y[53]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron54_1
  function_36 neuron54_1 (
      .a(input_layer[978]),
      .b(input_layer[603]),
      .c(input_layer[191]),
      .d(input_layer[1498]),
      .e(input_layer[287]),
      .f(~input_layer[878]),
      .y(Y[54]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron55_1
  function_37 neuron55_1 (
      .a(input_layer[1039]),
      .b(input_layer[1494]),
      .c(input_layer[159]),
      .d(~input_layer[628]),
      .e(~input_layer[1087]),
      .f(input_layer[1556]),
      .y(Y[55]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron56_1
  function_27 neuron56_1 (
      .a(~input_layer[1134]),
      .b(input_layer[907]),
      .c(~input_layer[517]),
      .y(Y[56]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_38 for neuron57_1
  function_38 neuron57_1 (
      .a(~input_layer[718]),
      .b(input_layer[1539]),
      .c(~input_layer[422]),
      .d(~input_layer[589]),
      .e(~input_layer[792]),
      .f(~input_layer[910]),
      .y(Y[57]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron58_1
  function_39 neuron58_1 (
      .a(input_layer[1026]),
      .b(~input_layer[1355]),
      .c(input_layer[525]),
      .y(Y[58]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron59_1
  function_40 neuron59_1 (
      .a(input_layer[1054]),
      .b(input_layer[1165]),
      .c(input_layer[312]),
      .d(~input_layer[821]),
      .e(input_layer[1197]),
      .f(input_layer[773]),
      .y(Y[59]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron60_1
  function_29 neuron60_1 (
      .a(~input_layer[1190]),
      .b(~input_layer[916]),
      .y(Y[60]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_41 for neuron61_1
  function_41 neuron61_1 (
      .a(input_layer[315]),
      .b(input_layer[372]),
      .c(~input_layer[1255]),
      .d(input_layer[940]),
      .e(input_layer[902]),
      .y(Y[61]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron62_1
  function_16 neuron62_1 (
      .a(input_layer[1358]),
      .b(~input_layer[364]),
      .y(Y[62]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron63_1
  function_4 neuron63_1 (
      .a(~input_layer[1027]),
      .b(input_layer[534]),
      .c(input_layer[530]),
      .d(~input_layer[1378]),
      .e(~input_layer[441]),
      .y(Y[63]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron64_1
  function_42 neuron64_1 (
      .a(input_layer[1126]),
      .b(input_layer[197]),
      .c(~input_layer[752]),
      .d(input_layer[1293]),
      .y(Y[64]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron65_1
  function_43 neuron65_1 (
      .a(~input_layer[1370]),
      .b(input_layer[212]),
      .c(~input_layer[547]),
      .d(input_layer[1067]),
      .e(input_layer[1253]),
      .f(input_layer[1517]),
      .y(Y[65]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron66_1
  function_44 neuron66_1 (
      .a(~input_layer[692]),
      .b(~input_layer[1488]),
      .c(input_layer[1157]),
      .d(~input_layer[770]),
      .e(~input_layer[859]),
      .y(Y[66]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron67_1
  function_19 neuron67_1 (
      .a(~input_layer[435]),
      .b(~input_layer[681]),
      .c(input_layer[751]),
      .d(~input_layer[268]),
      .y(Y[67]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron68_1
  function_27 neuron68_1 (
      .a(~input_layer[1330]),
      .b(~input_layer[641]),
      .c(~input_layer[582]),
      .y(Y[68]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron69_1
  function_27 neuron69_1 (
      .a(~input_layer[513]),
      .b(~input_layer[1549]),
      .c(~input_layer[137]),
      .y(Y[69]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron70_1
  function_45 neuron70_1 (
      .a(input_layer[518]),
      .b(input_layer[1364]),
      .c(input_layer[827]),
      .d(~input_layer[352]),
      .e(input_layer[1309]),
      .f(input_layer[564]),
      .y(Y[70]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron71_1
  function_46 neuron71_1 (
      .a(input_layer[1140]),
      .b(input_layer[1423]),
      .c(input_layer[732]),
      .d(input_layer[504]),
      .e(input_layer[1174]),
      .y(Y[71]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron72_1
  function_47 neuron72_1 (
      .a(input_layer[520]),
      .b(input_layer[1166]),
      .c(input_layer[770]),
      .d(input_layer[793]),
      .e(input_layer[653]),
      .y(Y[72]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron73_1
  function_48 neuron73_1 (
      .a(input_layer[1016]),
      .b(input_layer[304]),
      .c(input_layer[779]),
      .d(~input_layer[268]),
      .e(input_layer[1014]),
      .y(Y[73]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron74_1
  function_31 neuron74_1 (
      .a(~input_layer[1320]),
      .b(input_layer[1540]),
      .c(~input_layer[549]),
      .d(input_layer[352]),
      .y(Y[74]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron75_1
  function_49 neuron75_1 (
      .a(input_layer[585]),
      .b(~input_layer[544]),
      .c(input_layer[1160]),
      .d(~input_layer[1295]),
      .e(~input_layer[217]),
      .y(Y[75]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron76_1
  function_24 neuron76_1 (
      .a(input_layer[481]),
      .b(~input_layer[900]),
      .c(~input_layer[1295]),
      .y(Y[76]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron77_1
  function_16 neuron77_1 (
      .a(input_layer[637]),
      .b(input_layer[661]),
      .y(Y[77]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_41 for neuron78_1
  function_41 neuron78_1 (
      .a(input_layer[1021]),
      .b(input_layer[992]),
      .c(~input_layer[686]),
      .d(input_layer[1153]),
      .e(input_layer[503]),
      .y(Y[78]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron79_1
  function_48 neuron79_1 (
      .a(input_layer[878]),
      .b(input_layer[1181]),
      .c(input_layer[1168]),
      .d(input_layer[1363]),
      .e(input_layer[502]),
      .y(Y[79]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron80_1
  function_17 neuron80_1 (
      .a(input_layer[1053]),
      .b(input_layer[936]),
      .c(input_layer[403]),
      .y(Y[80]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron81_1
  function_39 neuron81_1 (
      .a(input_layer[606]),
      .b(input_layer[700]),
      .c(~input_layer[735]),
      .y(Y[81]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron82_1
  function_8 neuron82_1 (
      .a(input_layer[928]),
      .b(input_layer[1541]),
      .c(input_layer[563]),
      .d(input_layer[911]),
      .y(Y[82]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron83_1
  function_30 neuron83_1 (
      .a(~input_layer[1135]),
      .b(~input_layer[1307]),
      .c(~input_layer[1443]),
      .d(input_layer[1419]),
      .y(Y[83]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[84] = 1'b0;

  // instantiate function_50 for neuron85_1
  function_50 neuron85_1 (
      .a(~input_layer[869]),
      .b(input_layer[1327]),
      .c(input_layer[1242]),
      .d(~input_layer[1341]),
      .e(input_layer[25]),
      .f(~input_layer[0]),
      .y(Y[85]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron86_1
  function_3 neuron86_1 (
      .a(~input_layer[1383]),
      .b(~input_layer[1475]),
      .c(input_layer[1098]),
      .d(~input_layer[494]),
      .y(Y[86]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron87_1
  function_8 neuron87_1 (
      .a(input_layer[926]),
      .b(input_layer[131]),
      .c(~input_layer[968]),
      .d(~input_layer[434]),
      .y(Y[87]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_51 for neuron88_1
  function_51 neuron88_1 (
      .a(input_layer[1032]),
      .b(~input_layer[1132]),
      .c(~input_layer[800]),
      .d(~input_layer[525]),
      .e(input_layer[899]),
      .f(input_layer[27]),
      .y(Y[88]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron89_1
  function_52 neuron89_1 (
      .a(~input_layer[1202]),
      .b(input_layer[1474]),
      .c(~input_layer[501]),
      .d(input_layer[1338]),
      .e(~input_layer[64]),
      .f(~input_layer[1399]),
      .y(Y[89]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron90_1
  function_19 neuron90_1 (
      .a(~input_layer[1171]),
      .b(~input_layer[508]),
      .c(input_layer[391]),
      .d(input_layer[1254]),
      .y(Y[90]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron91_1
  function_8 neuron91_1 (
      .a(~input_layer[1256]),
      .b(input_layer[948]),
      .c(input_layer[1273]),
      .d(~input_layer[549]),
      .y(Y[91]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron92_1
  function_0 neuron92_1 (
      .a(input_layer[94]),
      .b(~input_layer[1033]),
      .c(~input_layer[962]),
      .d(~input_layer[116]),
      .e(~input_layer[1010]),
      .y(Y[92]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron93_1
  function_3 neuron93_1 (
      .a(~input_layer[1481]),
      .b(~input_layer[148]),
      .c(~input_layer[196]),
      .d(input_layer[318]),
      .y(Y[93]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron94_1
  function_53 neuron94_1 (
      .a(input_layer[1021]),
      .b(input_layer[184]),
      .c(input_layer[461]),
      .d(~input_layer[93]),
      .e(~input_layer[1532]),
      .f(~input_layer[725]),
      .y(Y[94]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron95_1
  function_3 neuron95_1 (
      .a(~input_layer[1081]),
      .b(~input_layer[323]),
      .c(~input_layer[934]),
      .d(input_layer[861]),
      .y(Y[95]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron96_1
  function_29 neuron96_1 (
      .a(~input_layer[1182]),
      .b(input_layer[579]),
      .y(Y[96]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron97_1
  function_54 neuron97_1 (
      .a(input_layer[440]),
      .b(~input_layer[793]),
      .c(input_layer[178]),
      .d(input_layer[1372]),
      .e(~input_layer[616]),
      .f(input_layer[121]),
      .y(Y[97]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron98_1
  function_55 neuron98_1 (
      .a(~input_layer[804]),
      .b(~input_layer[996]),
      .c(input_layer[520]),
      .d(~input_layer[889]),
      .e(~input_layer[1043]),
      .y(Y[98]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron99_1
  function_56 neuron99_1 (
      .a(input_layer[557]),
      .b(~input_layer[969]),
      .c(~input_layer[218]),
      .d(~input_layer[366]),
      .e(input_layer[1082]),
      .y(Y[99]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron100_1
  function_57 neuron100_1 (
      .a(input_layer[476]),
      .b(input_layer[418]),
      .c(~input_layer[437]),
      .d(~input_layer[795]),
      .e(input_layer[1465]),
      .f(input_layer[335]),
      .y(Y[100]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron101_1
  function_42 neuron101_1 (
      .a(input_layer[1429]),
      .b(input_layer[1466]),
      .c(input_layer[1381]),
      .d(input_layer[73]),
      .y(Y[101]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron102_1
  function_19 neuron102_1 (
      .a(~input_layer[689]),
      .b(~input_layer[638]),
      .c(input_layer[1035]),
      .d(~input_layer[217]),
      .y(Y[102]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron103_1
  function_16 neuron103_1 (
      .a(~input_layer[810]),
      .b(input_layer[1490]),
      .y(Y[103]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron104_1
  function_42 neuron104_1 (
      .a(input_layer[296]),
      .b(input_layer[271]),
      .c(input_layer[1111]),
      .d(~input_layer[1425]),
      .y(Y[104]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_58 for neuron105_1
  function_58 neuron105_1 (
      .a(input_layer[774]),
      .b(~input_layer[702]),
      .c(input_layer[1168]),
      .d(~input_layer[1322]),
      .e(input_layer[248]),
      .f(input_layer[1198]),
      .y(Y[105]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron106_1
  function_59 neuron106_1 (
      .a(input_layer[1248]),
      .b(input_layer[1187]),
      .c(input_layer[1548]),
      .d(input_layer[757]),
      .e(input_layer[993]),
      .f(~input_layer[1526]),
      .y(Y[106]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron107_1
  function_42 neuron107_1 (
      .a(input_layer[291]),
      .b(input_layer[452]),
      .c(input_layer[1152]),
      .d(input_layer[176]),
      .y(Y[107]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron108_1
  function_60 neuron108_1 (
      .a(input_layer[1492]),
      .b(~input_layer[432]),
      .c(input_layer[1546]),
      .d(~input_layer[1213]),
      .e(input_layer[839]),
      .y(Y[108]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron109_1
  function_0 neuron109_1 (
      .a(~input_layer[1429]),
      .b(~input_layer[1487]),
      .c(~input_layer[544]),
      .d(~input_layer[618]),
      .e(~input_layer[374]),
      .y(Y[109]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron110_1
  function_39 neuron110_1 (
      .a(input_layer[698]),
      .b(input_layer[666]),
      .c(~input_layer[892]),
      .y(Y[110]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron111_1
  function_39 neuron111_1 (
      .a(~input_layer[1053]),
      .b(input_layer[768]),
      .c(input_layer[83]),
      .y(Y[111]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron112_1
  function_29 neuron112_1 (
      .a(~input_layer[1266]),
      .b(input_layer[767]),
      .y(Y[112]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron113_1
  function_21 neuron113_1 (
      .a(input_layer[1330]),
      .b(~input_layer[513]),
      .c(~input_layer[1365]),
      .d(input_layer[1188]),
      .e(input_layer[275]),
      .y(Y[113]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron114_1
  function_0 neuron114_1 (
      .a(~input_layer[453]),
      .b(~input_layer[1086]),
      .c(~input_layer[232]),
      .d(~input_layer[1204]),
      .e(input_layer[415]),
      .y(Y[114]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron115_1
  function_61 neuron115_1 (
      .a(~input_layer[978]),
      .b(~input_layer[213]),
      .c(input_layer[1308]),
      .d(input_layer[1298]),
      .e(~input_layer[307]),
      .f(input_layer[939]),
      .y(Y[115]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron116_1
  function_7 neuron116_1 (
      .a(input_layer[919]),
      .b(input_layer[700]),
      .c(~input_layer[545]),
      .d(~input_layer[854]),
      .y(Y[116]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron117_1
  function_12 neuron117_1 (
      .a(input_layer[1136]),
      .b(~input_layer[804]),
      .c(~input_layer[1301]),
      .y(Y[117]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron118_1
  function_62 neuron118_1 (
      .a(input_layer[1023]),
      .b(input_layer[1442]),
      .c(~input_layer[646]),
      .d(input_layer[350]),
      .e(input_layer[1200]),
      .f(input_layer[389]),
      .y(Y[118]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron119_1
  function_27 neuron119_1 (
      .a(~input_layer[1070]),
      .b(~input_layer[1544]),
      .c(~input_layer[944]),
      .y(Y[119]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron120_1
  function_40 neuron120_1 (
      .a(input_layer[398]),
      .b(input_layer[834]),
      .c(~input_layer[1248]),
      .d(input_layer[1281]),
      .e(~input_layer[1210]),
      .f(~input_layer[417]),
      .y(Y[120]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron121_1
  function_3 neuron121_1 (
      .a(~input_layer[882]),
      .b(~input_layer[1129]),
      .c(~input_layer[423]),
      .d(~input_layer[1010]),
      .y(Y[121]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron122_1
  function_3 neuron122_1 (
      .a(~input_layer[861]),
      .b(~input_layer[1471]),
      .c(~input_layer[801]),
      .d(~input_layer[398]),
      .y(Y[122]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron123_1
  function_14 neuron123_1 (
      .a(input_layer[1478]),
      .b(~input_layer[1030]),
      .c(input_layer[1246]),
      .d(input_layer[1380]),
      .e(~input_layer[121]),
      .f(input_layer[606]),
      .y(Y[123]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron124_1
  function_63 neuron124_1 (
      .a(~input_layer[876]),
      .b(input_layer[551]),
      .c(input_layer[669]),
      .d(input_layer[373]),
      .e(input_layer[415]),
      .y(Y[124]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron125_1
  function_26 neuron125_1 (
      .a(input_layer[800]),
      .y(Y[125]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron126_1
  function_29 neuron126_1 (
      .a(~input_layer[739]),
      .b(input_layer[461]),
      .y(Y[126]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[127] = 1'b0;

  // instantiate function_64 for neuron128_1
  function_64 neuron128_1 (
      .a(input_layer[721]),
      .b(~input_layer[1416]),
      .c(input_layer[307]),
      .d(input_layer[1090]),
      .e(~input_layer[855]),
      .y(Y[128]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron129_1
  function_65 neuron129_1 (
      .a(~input_layer[603]),
      .b(~input_layer[641]),
      .c(input_layer[904]),
      .d(input_layer[1222]),
      .e(input_layer[154]),
      .f(~input_layer[121]),
      .y(Y[129]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron130_1
  function_57 neuron130_1 (
      .a(input_layer[411]),
      .b(input_layer[1311]),
      .c(~input_layer[822]),
      .d(~input_layer[1334]),
      .e(input_layer[722]),
      .f(~input_layer[116]),
      .y(Y[130]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_66 for neuron131_1
  function_66 neuron131_1 (
      .a(input_layer[966]),
      .b(~input_layer[755]),
      .c(~input_layer[603]),
      .d(~input_layer[646]),
      .e(~input_layer[1557]),
      .f(~input_layer[846]),
      .y(Y[131]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron132_1
  function_1 neuron132_1 (
      .a(~input_layer[1137]),
      .b(input_layer[823]),
      .c(~input_layer[1136]),
      .d(~input_layer[413]),
      .y(Y[132]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron133_1
  function_17 neuron133_1 (
      .a(input_layer[947]),
      .b(input_layer[1278]),
      .c(~input_layer[930]),
      .y(Y[133]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron134_1
  function_42 neuron134_1 (
      .a(input_layer[914]),
      .b(input_layer[903]),
      .c(input_layer[1335]),
      .d(input_layer[1389]),
      .y(Y[134]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron135_1
  function_67 neuron135_1 (
      .a(~input_layer[1137]),
      .b(~input_layer[1195]),
      .c(~input_layer[509]),
      .d(~input_layer[1362]),
      .e(~input_layer[1171]),
      .y(Y[135]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron136_1
  function_0 neuron136_1 (
      .a(~input_layer[437]),
      .b(input_layer[1387]),
      .c(~input_layer[1074]),
      .d(~input_layer[93]),
      .e(~input_layer[727]),
      .y(Y[136]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron137_1
  function_7 neuron137_1 (
      .a(~input_layer[637]),
      .b(input_layer[1117]),
      .c(input_layer[869]),
      .d(input_layer[274]),
      .y(Y[137]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron138_1
  function_8 neuron138_1 (
      .a(input_layer[964]),
      .b(~input_layer[1369]),
      .c(input_layer[76]),
      .d(input_layer[479]),
      .y(Y[138]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_68 for neuron139_1
  function_68 neuron139_1 (
      .a(input_layer[753]),
      .b(~input_layer[1439]),
      .c(~input_layer[848]),
      .d(input_layer[314]),
      .e(~input_layer[616]),
      .f(input_layer[339]),
      .y(Y[139]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron140_1
  function_4 neuron140_1 (
      .a(~input_layer[409]),
      .b(input_layer[754]),
      .c(~input_layer[1046]),
      .d(~input_layer[847]),
      .e(input_layer[121]),
      .y(Y[140]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron141_1
  function_37 neuron141_1 (
      .a(input_layer[194]),
      .b(input_layer[240]),
      .c(~input_layer[611]),
      .d(~input_layer[602]),
      .e(input_layer[127]),
      .f(input_layer[518]),
      .y(Y[141]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron142_1
  function_69 neuron142_1 (
      .a(input_layer[444]),
      .b(~input_layer[749]),
      .c(~input_layer[995]),
      .d(~input_layer[832]),
      .e(input_layer[902]),
      .f(~input_layer[23]),
      .y(Y[142]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron143_1
  function_70 neuron143_1 (
      .a(~input_layer[1023]),
      .b(input_layer[1307]),
      .c(~input_layer[890]),
      .d(input_layer[308]),
      .e(input_layer[68]),
      .f(input_layer[25]),
      .y(Y[143]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_71 for neuron144_1
  function_71 neuron144_1 (
      .a(input_layer[875]),
      .b(~input_layer[486]),
      .c(input_layer[932]),
      .d(input_layer[1530]),
      .e(input_layer[289]),
      .f(input_layer[1448]),
      .y(Y[144]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron145_1
  function_12 neuron145_1 (
      .a(input_layer[268]),
      .b(input_layer[302]),
      .c(~input_layer[1358]),
      .y(Y[145]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron146_1
  function_29 neuron146_1 (
      .a(~input_layer[1240]),
      .b(~input_layer[478]),
      .y(Y[146]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron147_1
  function_46 neuron147_1 (
      .a(~input_layer[752]),
      .b(input_layer[850]),
      .c(input_layer[1003]),
      .d(input_layer[470]),
      .e(~input_layer[702]),
      .y(Y[147]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron148_1
  function_29 neuron148_1 (
      .a(input_layer[552]),
      .b(~input_layer[741]),
      .y(Y[148]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron149_1
  function_72 neuron149_1 (
      .a(input_layer[1431]),
      .b(input_layer[1424]),
      .c(~input_layer[260]),
      .d(~input_layer[611]),
      .e(input_layer[560]),
      .y(Y[149]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_73 for neuron150_1
  function_73 neuron150_1 (
      .a(~input_layer[1383]),
      .b(input_layer[1219]),
      .c(input_layer[463]),
      .d(input_layer[780]),
      .e(~input_layer[169]),
      .f(~input_layer[133]),
      .y(Y[150]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron151_1
  function_74 neuron151_1 (
      .a(~input_layer[1249]),
      .b(~input_layer[512]),
      .c(~input_layer[1192]),
      .d(~input_layer[1409]),
      .e(input_layer[1448]),
      .f(~input_layer[28]),
      .y(Y[151]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron152_1
  function_75 neuron152_1 (
      .a(input_layer[600]),
      .b(~input_layer[330]),
      .c(input_layer[419]),
      .d(~input_layer[315]),
      .e(~input_layer[978]),
      .y(Y[152]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron153_1
  function_76 neuron153_1 (
      .a(input_layer[406]),
      .b(input_layer[611]),
      .c(input_layer[181]),
      .d(input_layer[562]),
      .e(~input_layer[909]),
      .f(input_layer[122]),
      .y(Y[153]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_77 for neuron154_1
  function_77 neuron154_1 (
      .a(input_layer[803]),
      .b(~input_layer[307]),
      .c(input_layer[620]),
      .d(~input_layer[254]),
      .e(input_layer[1207]),
      .f(input_layer[333]),
      .y(Y[154]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron155_1
  function_45 neuron155_1 (
      .a(input_layer[572]),
      .b(input_layer[1491]),
      .c(~input_layer[364]),
      .d(input_layer[124]),
      .e(~input_layer[350]),
      .f(input_layer[317]),
      .y(Y[155]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron156_1
  function_17 neuron156_1 (
      .a(input_layer[762]),
      .b(input_layer[993]),
      .c(input_layer[296]),
      .y(Y[156]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron157_1
  function_78 neuron157_1 (
      .a(~input_layer[751]),
      .b(~input_layer[608]),
      .c(~input_layer[134]),
      .d(~input_layer[1446]),
      .e(~input_layer[1182]),
      .f(~input_layer[420]),
      .y(Y[157]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron158_1
  function_27 neuron158_1 (
      .a(~input_layer[1056]),
      .b(~input_layer[1201]),
      .c(input_layer[741]),
      .y(Y[158]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_79 for neuron159_1
  function_79 neuron159_1 (
      .a(~input_layer[934]),
      .b(~input_layer[589]),
      .c(input_layer[193]),
      .d(~input_layer[78]),
      .e(~input_layer[129]),
      .f(input_layer[1241]),
      .y(Y[159]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_80 for neuron160_1
  function_80 neuron160_1 (
      .a(input_layer[578]),
      .b(~input_layer[1154]),
      .c(~input_layer[1237]),
      .d(~input_layer[1270]),
      .e(~input_layer[1189]),
      .f(~input_layer[1329]),
      .y(Y[160]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_81 for neuron161_1
  function_81 neuron161_1 (
      .a(input_layer[360]),
      .b(~input_layer[978]),
      .c(input_layer[1020]),
      .d(input_layer[274]),
      .e(~input_layer[704]),
      .f(input_layer[540]),
      .y(Y[161]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron162_1
  function_82 neuron162_1 (
      .a(~input_layer[651]),
      .b(input_layer[810]),
      .c(~input_layer[423]),
      .d(input_layer[1198]),
      .e(~input_layer[1556]),
      .f(input_layer[901]),
      .y(Y[162]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron163_1
  function_27 neuron163_1 (
      .a(~input_layer[1313]),
      .b(~input_layer[1275]),
      .c(input_layer[1148]),
      .y(Y[163]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_83 for neuron164_1
  function_83 neuron164_1 (
      .a(input_layer[1479]),
      .b(~input_layer[908]),
      .c(~input_layer[415]),
      .d(~input_layer[1307]),
      .e(~input_layer[129]),
      .y(Y[164]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron165_1
  function_17 neuron165_1 (
      .a(input_layer[918]),
      .b(input_layer[869]),
      .c(input_layer[184]),
      .y(Y[165]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron166_1
  function_84 neuron166_1 (
      .a(~input_layer[324]),
      .b(~input_layer[878]),
      .c(input_layer[1035]),
      .d(input_layer[536]),
      .e(input_layer[392]),
      .y(Y[166]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron167_1
  function_85 neuron167_1 (
      .a(input_layer[1039]),
      .b(~input_layer[1155]),
      .c(input_layer[830]),
      .d(input_layer[469]),
      .e(input_layer[1009]),
      .f(input_layer[24]),
      .y(Y[167]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron168_1
  function_45 neuron168_1 (
      .a(input_layer[198]),
      .b(~input_layer[857]),
      .c(input_layer[252]),
      .d(input_layer[1501]),
      .e(input_layer[1199]),
      .f(input_layer[99]),
      .y(Y[168]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron169_1
  function_24 neuron169_1 (
      .a(~input_layer[1150]),
      .b(~input_layer[386]),
      .c(input_layer[1333]),
      .y(Y[169]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron170_1
  function_26 neuron170_1 (
      .a(input_layer[633]),
      .y(Y[170]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron171_1
  function_27 neuron171_1 (
      .a(~input_layer[1494]),
      .b(input_layer[976]),
      .c(~input_layer[1413]),
      .y(Y[171]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron172_1
  function_16 neuron172_1 (
      .a(input_layer[823]),
      .b(input_layer[820]),
      .y(Y[172]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_86 for neuron173_1
  function_86 neuron173_1 (
      .a(input_layer[249]),
      .b(input_layer[1191]),
      .c(input_layer[1012]),
      .d(input_layer[1075]),
      .e(~input_layer[1041]),
      .f(~input_layer[203]),
      .y(Y[173]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron174_1
  function_47 neuron174_1 (
      .a(input_layer[1368]),
      .b(input_layer[1421]),
      .c(input_layer[345]),
      .d(input_layer[789]),
      .e(input_layer[755]),
      .y(Y[174]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron175_1
  function_56 neuron175_1 (
      .a(input_layer[716]),
      .b(~input_layer[498]),
      .c(input_layer[1470]),
      .d(~input_layer[432]),
      .e(~input_layer[1272]),
      .y(Y[175]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron176_1
  function_87 neuron176_1 (
      .a(input_layer[1333]),
      .b(~input_layer[1044]),
      .c(~input_layer[801]),
      .d(input_layer[304]),
      .e(input_layer[42]),
      .y(Y[176]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron177_1
  function_42 neuron177_1 (
      .a(input_layer[389]),
      .b(input_layer[1293]),
      .c(~input_layer[864]),
      .d(input_layer[615]),
      .y(Y[177]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron178_1
  function_27 neuron178_1 (
      .a(~input_layer[527]),
      .b(~input_layer[1078]),
      .c(~input_layer[1079]),
      .y(Y[178]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron179_1
  function_19 neuron179_1 (
      .a(~input_layer[485]),
      .b(~input_layer[832]),
      .c(input_layer[314]),
      .d(input_layer[333]),
      .y(Y[179]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_88 for neuron180_1
  function_88 neuron180_1 (
      .a(~input_layer[529]),
      .b(~input_layer[720]),
      .c(input_layer[25]),
      .d(input_layer[842]),
      .e(~input_layer[945]),
      .f(input_layer[64]),
      .y(Y[180]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron181_1
  function_89 neuron181_1 (
      .a(input_layer[1081]),
      .b(input_layer[1139]),
      .c(~input_layer[1125]),
      .d(~input_layer[381]),
      .e(~input_layer[674]),
      .y(Y[181]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron182_1
  function_40 neuron182_1 (
      .a(input_layer[198]),
      .b(~input_layer[858]),
      .c(input_layer[1156]),
      .d(input_layer[646]),
      .e(input_layer[272]),
      .f(input_layer[122]),
      .y(Y[182]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron183_1
  function_90 neuron183_1 (
      .a(~input_layer[256]),
      .b(input_layer[1426]),
      .c(~input_layer[361]),
      .d(input_layer[413]),
      .e(~input_layer[1030]),
      .y(Y[183]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron184_1
  function_91 neuron184_1 (
      .a(~input_layer[876]),
      .b(input_layer[1499]),
      .c(~input_layer[328]),
      .d(~input_layer[460]),
      .e(~input_layer[272]),
      .y(Y[184]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron185_1
  function_55 neuron185_1 (
      .a(~input_layer[404]),
      .b(~input_layer[554]),
      .c(~input_layer[1321]),
      .d(~input_layer[435]),
      .e(~input_layer[1216]),
      .y(Y[185]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron186_1
  function_92 neuron186_1 (
      .a(input_layer[1477]),
      .b(input_layer[1474]),
      .c(input_layer[454]),
      .d(input_layer[1084]),
      .e(~input_layer[231]),
      .f(~input_layer[1395]),
      .y(Y[186]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron187_1
  function_92 neuron187_1 (
      .a(input_layer[354]),
      .b(input_layer[1053]),
      .c(input_layer[1043]),
      .d(input_layer[90]),
      .e(~input_layer[981]),
      .f(input_layer[120]),
      .y(Y[187]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron188_1
  function_93 neuron188_1 (
      .a(~input_layer[200]),
      .b(input_layer[1437]),
      .c(input_layer[1445]),
      .d(~input_layer[1475]),
      .e(input_layer[331]),
      .y(Y[188]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron189_1
  function_12 neuron189_1 (
      .a(input_layer[695]),
      .b(input_layer[331]),
      .c(~input_layer[1499]),
      .y(Y[189]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron190_1
  function_24 neuron190_1 (
      .a(~input_layer[1142]),
      .b(~input_layer[217]),
      .c(~input_layer[913]),
      .y(Y[190]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron191_1
  function_12 neuron191_1 (
      .a(input_layer[379]),
      .b(input_layer[262]),
      .c(~input_layer[1169]),
      .y(Y[191]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron192_1
  function_3 neuron192_1 (
      .a(~input_layer[1434]),
      .b(~input_layer[927]),
      .c(~input_layer[330]),
      .d(input_layer[486]),
      .y(Y[192]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_94 for neuron193_1
  function_94 neuron193_1 (
      .a(input_layer[1110]),
      .b(~input_layer[415]),
      .c(input_layer[1109]),
      .d(input_layer[1106]),
      .e(~input_layer[15]),
      .f(input_layer[73]),
      .y(Y[193]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron194_1
  function_95 neuron194_1 (
      .a(input_layer[1544]),
      .b(~input_layer[1251]),
      .c(~input_layer[263]),
      .d(input_layer[83]),
      .y(Y[194]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron195_1
  function_96 neuron195_1 (
      .a(~input_layer[975]),
      .b(~input_layer[183]),
      .c(input_layer[665]),
      .d(input_layer[586]),
      .y(Y[195]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron196_1
  function_97 neuron196_1 (
      .a(~input_layer[512]),
      .b(~input_layer[465]),
      .c(~input_layer[398]),
      .d(input_layer[998]),
      .e(input_layer[310]),
      .y(Y[196]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron197_1
  function_27 neuron197_1 (
      .a(~input_layer[441]),
      .b(input_layer[699]),
      .c(~input_layer[585]),
      .y(Y[197]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_98 for neuron198_1
  function_98 neuron198_1 (
      .a(~input_layer[239]),
      .b(~input_layer[192]),
      .c(input_layer[910]),
      .d(input_layer[1143]),
      .e(~input_layer[1368]),
      .f(input_layer[430]),
      .y(Y[198]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron199_1
  function_8 neuron199_1 (
      .a(input_layer[208]),
      .b(input_layer[237]),
      .c(~input_layer[1133]),
      .d(input_layer[264]),
      .y(Y[199]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron200_1
  function_99 neuron200_1 (
      .a(input_layer[1486]),
      .b(~input_layer[991]),
      .c(input_layer[572]),
      .d(~input_layer[817]),
      .e(~input_layer[1095]),
      .y(Y[200]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron201_1
  function_8 neuron201_1 (
      .a(input_layer[1331]),
      .b(input_layer[946]),
      .c(input_layer[949]),
      .d(~input_layer[686]),
      .y(Y[201]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron202_1
  function_100 neuron202_1 (
      .a(~input_layer[608]),
      .b(~input_layer[700]),
      .c(input_layer[525]),
      .d(input_layer[1435]),
      .e(~input_layer[1438]),
      .f(~input_layer[233]),
      .y(Y[202]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_101 for neuron203_1
  function_101 neuron203_1 (
      .a(input_layer[921]),
      .b(~input_layer[1408]),
      .c(input_layer[926]),
      .d(input_layer[159]),
      .e(~input_layer[443]),
      .f(~input_layer[557]),
      .y(Y[203]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron204_1
  function_29 neuron204_1 (
      .a(~input_layer[555]),
      .b(input_layer[964]),
      .y(Y[204]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron205_1
  function_74 neuron205_1 (
      .a(~input_layer[767]),
      .b(~input_layer[575]),
      .c(~input_layer[1022]),
      .d(~input_layer[1155]),
      .e(~input_layer[948]),
      .f(input_layer[1458]),
      .y(Y[205]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_102 for neuron206_1
  function_102 neuron206_1 (
      .a(~input_layer[301]),
      .b(~input_layer[1236]),
      .c(~input_layer[1268]),
      .d(input_layer[769]),
      .e(input_layer[424]),
      .f(input_layer[22]),
      .y(Y[206]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron207_1
  function_27 neuron207_1 (
      .a(~input_layer[599]),
      .b(~input_layer[945]),
      .c(input_layer[526]),
      .y(Y[207]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron208_1
  function_29 neuron208_1 (
      .a(~input_layer[384]),
      .b(input_layer[1088]),
      .y(Y[208]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron209_1
  function_72 neuron209_1 (
      .a(~input_layer[88]),
      .b(~input_layer[1079]),
      .c(input_layer[235]),
      .d(input_layer[374]),
      .e(input_layer[493]),
      .y(Y[209]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_103 for neuron210_1
  function_103 neuron210_1 (
      .a(~input_layer[1422]),
      .b(input_layer[421]),
      .c(input_layer[551]),
      .d(input_layer[158]),
      .e(input_layer[73]),
      .f(~input_layer[111]),
      .y(Y[210]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron211_1
  function_104 neuron211_1 (
      .a(input_layer[296]),
      .b(input_layer[1273]),
      .c(input_layer[373]),
      .d(~input_layer[1013]),
      .e(~input_layer[56]),
      .f(~input_layer[281]),
      .y(Y[211]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_105 for neuron212_1
  function_105 neuron212_1 (
      .a(~input_layer[328]),
      .b(~input_layer[583]),
      .c(input_layer[1127]),
      .d(input_layer[476]),
      .e(input_layer[891]),
      .y(Y[212]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron213_1
  function_3 neuron213_1 (
      .a(~input_layer[537]),
      .b(~input_layer[243]),
      .c(~input_layer[891]),
      .d(input_layer[1195]),
      .y(Y[213]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron214_1
  function_11 neuron214_1 (
      .a(input_layer[803]),
      .b(~input_layer[1547]),
      .c(~input_layer[234]),
      .d(~input_layer[707]),
      .y(Y[214]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron215_1
  function_106 neuron215_1 (
      .a(input_layer[1427]),
      .b(~input_layer[445]),
      .c(input_layer[1415]),
      .d(input_layer[685]),
      .y(Y[215]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron216_1
  function_107 neuron216_1 (
      .a(~input_layer[1198]),
      .b(~input_layer[1527]),
      .c(input_layer[218]),
      .d(~input_layer[1223]),
      .e(input_layer[590]),
      .y(Y[216]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_108 for neuron217_1
  function_108 neuron217_1 (
      .a(input_layer[1070]),
      .b(~input_layer[654]),
      .c(input_layer[1245]),
      .d(input_layer[288]),
      .e(input_layer[960]),
      .f(~input_layer[79]),
      .y(Y[217]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_109 for neuron218_1
  function_109 neuron218_1 (
      .a(input_layer[296]),
      .b(~input_layer[775]),
      .c(~input_layer[272]),
      .d(input_layer[653]),
      .e(~input_layer[71]),
      .f(~input_layer[838]),
      .y(Y[218]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron219_1
  function_67 neuron219_1 (
      .a(~input_layer[1185]),
      .b(~input_layer[1272]),
      .c(~input_layer[425]),
      .d(~input_layer[1336]),
      .e(~input_layer[903]),
      .y(Y[219]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_110 for neuron220_1
  function_110 neuron220_1 (
      .a(input_layer[682]),
      .b(~input_layer[973]),
      .c(~input_layer[456]),
      .d(input_layer[1384]),
      .e(~input_layer[835]),
      .f(~input_layer[986]),
      .y(Y[220]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron221_1
  function_27 neuron221_1 (
      .a(~input_layer[1025]),
      .b(~input_layer[966]),
      .c(input_layer[1308]),
      .y(Y[221]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_111 for neuron222_1
  function_111 neuron222_1 (
      .a(input_layer[430]),
      .b(~input_layer[82]),
      .c(input_layer[357]),
      .d(input_layer[355]),
      .e(input_layer[1295]),
      .y(Y[222]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron223_1
  function_100 neuron223_1 (
      .a(~input_layer[1141]),
      .b(~input_layer[945]),
      .c(input_layer[466]),
      .d(~input_layer[679]),
      .e(~input_layer[674]),
      .f(~input_layer[1024]),
      .y(Y[223]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron224_1
  function_27 neuron224_1 (
      .a(~input_layer[455]),
      .b(~input_layer[835]),
      .c(input_layer[980]),
      .y(Y[224]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron225_1
  function_29 neuron225_1 (
      .a(input_layer[366]),
      .b(~input_layer[1051]),
      .y(Y[225]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron226_1
  function_112 neuron226_1 (
      .a(~input_layer[699]),
      .b(~input_layer[390]),
      .c(input_layer[351]),
      .d(input_layer[655]),
      .e(input_layer[30]),
      .f(~input_layer[1563]),
      .y(Y[226]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron227_1
  function_113 neuron227_1 (
      .a(~input_layer[1191]),
      .b(input_layer[776]),
      .c(input_layer[131]),
      .d(~input_layer[1413]),
      .e(input_layer[507]),
      .y(Y[227]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_114 for neuron228_1
  function_114 neuron228_1 (
      .a(~input_layer[647]),
      .b(~input_layer[923]),
      .c(input_layer[1069]),
      .d(input_layer[755]),
      .e(~input_layer[1319]),
      .f(~input_layer[394]),
      .y(Y[228]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron229_1
  function_19 neuron229_1 (
      .a(~input_layer[1071]),
      .b(~input_layer[1353]),
      .c(~input_layer[1030]),
      .d(input_layer[792]),
      .y(Y[229]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron230_1
  function_99 neuron230_1 (
      .a(input_layer[359]),
      .b(input_layer[1024]),
      .c(~input_layer[1354]),
      .d(~input_layer[528]),
      .e(input_layer[1283]),
      .y(Y[230]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron231_1
  function_26 neuron231_1 (
      .a(~input_layer[1094]),
      .y(Y[231]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron232_1
  function_16 neuron232_1 (
      .a(input_layer[303]),
      .b(input_layer[1220]),
      .y(Y[232]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron233_1
  function_115 neuron233_1 (
      .a(~input_layer[1020]),
      .b(input_layer[1421]),
      .c(input_layer[517]),
      .d(~input_layer[77]),
      .e(input_layer[562]),
      .f(input_layer[489]),
      .y(Y[233]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron234_1
  function_42 neuron234_1 (
      .a(input_layer[919]),
      .b(input_layer[1238]),
      .c(input_layer[1113]),
      .d(~input_layer[981]),
      .y(Y[234]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron235_1
  function_116 neuron235_1 (
      .a(input_layer[973]),
      .b(~input_layer[1418]),
      .c(~input_layer[810]),
      .d(~input_layer[295]),
      .e(~input_layer[1211]),
      .f(~input_layer[84]),
      .y(Y[235]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron236_1
  function_117 neuron236_1 (
      .a(~input_layer[437]),
      .b(input_layer[1106]),
      .c(~input_layer[1383]),
      .d(input_layer[622]),
      .e(input_layer[1349]),
      .f(~input_layer[1286]),
      .y(Y[236]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_118 for neuron237_1
  function_118 neuron237_1 (
      .a(input_layer[540]),
      .b(~input_layer[266]),
      .c(input_layer[734]),
      .d(input_layer[1306]),
      .e(input_layer[654]),
      .f(~input_layer[248]),
      .y(Y[237]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron238_1
  function_119 neuron238_1 (
      .a(~input_layer[1029]),
      .b(~input_layer[714]),
      .c(~input_layer[548]),
      .d(~input_layer[907]),
      .e(input_layer[1066]),
      .y(Y[238]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron239_1
  function_18 neuron239_1 (
      .a(~input_layer[145]),
      .b(input_layer[1296]),
      .c(input_layer[876]),
      .d(~input_layer[775]),
      .e(input_layer[18]),
      .y(Y[239]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron240_1
  function_42 neuron240_1 (
      .a(input_layer[410]),
      .b(input_layer[552]),
      .c(input_layer[696]),
      .d(input_layer[1105]),
      .y(Y[240]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron241_1
  function_120 neuron241_1 (
      .a(input_layer[327]),
      .b(~input_layer[1482]),
      .c(input_layer[959]),
      .d(~input_layer[793]),
      .e(~input_layer[769]),
      .y(Y[241]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron242_1
  function_70 neuron242_1 (
      .a(~input_layer[534]),
      .b(input_layer[650]),
      .c(~input_layer[1466]),
      .d(~input_layer[1154]),
      .e(input_layer[216]),
      .f(~input_layer[1030]),
      .y(Y[242]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron243_1
  function_121 neuron243_1 (
      .a(input_layer[1133]),
      .b(input_layer[1220]),
      .c(~input_layer[159]),
      .d(input_layer[618]),
      .e(~input_layer[1420]),
      .y(Y[243]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_122 for neuron244_1
  function_122 neuron244_1 (
      .a(input_layer[909]),
      .b(~input_layer[306]),
      .c(~input_layer[1379]),
      .d(input_layer[913]),
      .e(input_layer[1341]),
      .f(input_layer[899]),
      .y(Y[244]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron245_1
  function_36 neuron245_1 (
      .a(input_layer[1414]),
      .b(input_layer[566]),
      .c(~input_layer[923]),
      .d(input_layer[1095]),
      .e(input_layer[734]),
      .f(input_layer[992]),
      .y(Y[245]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron246_1
  function_7 neuron246_1 (
      .a(input_layer[598]),
      .b(~input_layer[1368]),
      .c(input_layer[1180]),
      .d(input_layer[761]),
      .y(Y[246]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron247_1
  function_47 neuron247_1 (
      .a(input_layer[241]),
      .b(input_layer[554]),
      .c(input_layer[1212]),
      .d(input_layer[332]),
      .e(~input_layer[516]),
      .y(Y[247]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron248_1
  function_123 neuron248_1 (
      .a(input_layer[970]),
      .b(~input_layer[703]),
      .c(input_layer[1228]),
      .d(~input_layer[412]),
      .y(Y[248]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron249_1
  function_11 neuron249_1 (
      .a(~input_layer[870]),
      .b(~input_layer[333]),
      .c(input_layer[252]),
      .d(~input_layer[558]),
      .y(Y[249]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron250_1
  function_42 neuron250_1 (
      .a(input_layer[151]),
      .b(input_layer[941]),
      .c(input_layer[801]),
      .d(input_layer[1445]),
      .y(Y[250]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron251_1
  function_24 neuron251_1 (
      .a(~input_layer[689]),
      .b(input_layer[1146]),
      .c(~input_layer[1375]),
      .y(Y[251]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron252_1
  function_16 neuron252_1 (
      .a(input_layer[1297]),
      .b(~input_layer[1031]),
      .y(Y[252]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_124 for neuron253_1
  function_124 neuron253_1 (
      .a(~input_layer[325]),
      .b(~input_layer[196]),
      .c(input_layer[526]),
      .d(~input_layer[804]),
      .e(~input_layer[923]),
      .f(~input_layer[209]),
      .y(Y[253]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron254_1
  function_96 neuron254_1 (
      .a(~input_layer[1081]),
      .b(input_layer[822]),
      .c(~input_layer[1278]),
      .d(input_layer[1500]),
      .y(Y[254]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron255_1
  function_125 neuron255_1 (
      .a(input_layer[977]),
      .b(~input_layer[762]),
      .c(input_layer[601]),
      .d(~input_layer[861]),
      .e(input_layer[335]),
      .f(input_layer[56]),
      .y(Y[255]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron256_1
  function_29 neuron256_1 (
      .a(~input_layer[915]),
      .b(~input_layer[493]),
      .y(Y[256]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron257_1
  function_26 neuron257_1 (
      .a(input_layer[1310]),
      .y(Y[257]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron258_1
  function_17 neuron258_1 (
      .a(input_layer[762]),
      .b(input_layer[185]),
      .c(input_layer[1386]),
      .y(Y[258]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron259_1
  function_17 neuron259_1 (
      .a(input_layer[381]),
      .b(input_layer[1369]),
      .c(input_layer[1293]),
      .y(Y[259]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron260_1
  function_126 neuron260_1 (
      .a(~input_layer[371]),
      .b(~input_layer[1144]),
      .c(~input_layer[1129]),
      .d(~input_layer[946]),
      .e(input_layer[389]),
      .y(Y[260]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_127 for neuron261_1
  function_127 neuron261_1 (
      .a(input_layer[1414]),
      .b(~input_layer[821]),
      .c(input_layer[1303]),
      .d(input_layer[1154]),
      .e(input_layer[236]),
      .f(~input_layer[1013]),
      .y(Y[261]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron262_1
  function_128 neuron262_1 (
      .a(~input_layer[322]),
      .b(input_layer[1552]),
      .c(~input_layer[296]),
      .d(~input_layer[1095]),
      .y(Y[262]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron263_1
  function_100 neuron263_1 (
      .a(~input_layer[748]),
      .b(~input_layer[656]),
      .c(input_layer[866]),
      .d(~input_layer[1330]),
      .e(~input_layer[304]),
      .f(~input_layer[276]),
      .y(Y[263]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron264_1
  function_46 neuron264_1 (
      .a(input_layer[195]),
      .b(~input_layer[751]),
      .c(input_layer[1434]),
      .d(input_layer[531]),
      .e(input_layer[1145]),
      .y(Y[264]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron265_1
  function_8 neuron265_1 (
      .a(input_layer[414]),
      .b(input_layer[850]),
      .c(input_layer[951]),
      .d(input_layer[231]),
      .y(Y[265]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_129 for neuron266_1
  function_129 neuron266_1 (
      .a(input_layer[552]),
      .b(~input_layer[462]),
      .c(input_layer[1434]),
      .d(~input_layer[1514]),
      .e(input_layer[896]),
      .f(~input_layer[108]),
      .y(Y[266]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[267] = 1'b0;

  // instantiate function_130 for neuron268_1
  function_130 neuron268_1 (
      .a(~input_layer[1372]),
      .b(~input_layer[978]),
      .c(input_layer[419]),
      .d(~input_layer[669]),
      .e(input_layer[1163]),
      .f(~input_layer[724]),
      .y(Y[268]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_105 for neuron269_1
  function_105 neuron269_1 (
      .a(input_layer[636]),
      .b(~input_layer[1239]),
      .c(input_layer[584]),
      .d(input_layer[1132]),
      .e(~input_layer[1316]),
      .y(Y[269]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron270_1
  function_131 neuron270_1 (
      .a(~input_layer[774]),
      .b(input_layer[1375]),
      .c(~input_layer[915]),
      .d(input_layer[1359]),
      .e(~input_layer[210]),
      .f(input_layer[341]),
      .y(Y[270]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron271_1
  function_92 neuron271_1 (
      .a(input_layer[1485]),
      .b(input_layer[713]),
      .c(input_layer[321]),
      .d(input_layer[1437]),
      .e(input_layer[710]),
      .f(~input_layer[45]),
      .y(Y[271]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron272_1
  function_132 neuron272_1 (
      .a(input_layer[1077]),
      .b(input_layer[1252]),
      .c(~input_layer[140]),
      .d(input_layer[846]),
      .e(input_layer[405]),
      .f(~input_layer[1161]),
      .y(Y[272]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron273_1
  function_31 neuron273_1 (
      .a(~input_layer[1189]),
      .b(~input_layer[1263]),
      .c(input_layer[1470]),
      .d(input_layer[403]),
      .y(Y[273]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron274_1
  function_133 neuron274_1 (
      .a(~input_layer[1169]),
      .b(~input_layer[194]),
      .c(input_layer[620]),
      .d(input_layer[343]),
      .e(input_layer[487]),
      .f(~input_layer[1240]),
      .y(Y[274]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron275_1
  function_46 neuron275_1 (
      .a(input_layer[980]),
      .b(input_layer[648]),
      .c(input_layer[1069]),
      .d(~input_layer[367]),
      .e(input_layer[1557]),
      .y(Y[275]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron276_1
  function_26 neuron276_1 (
      .a(input_layer[533]),
      .y(Y[276]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron277_1
  function_17 neuron277_1 (
      .a(input_layer[1468]),
      .b(input_layer[1320]),
      .c(~input_layer[251]),
      .y(Y[277]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron278_1
  function_30 neuron278_1 (
      .a(~input_layer[927]),
      .b(input_layer[808]),
      .c(input_layer[354]),
      .d(input_layer[721]),
      .y(Y[278]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron279_1
  function_46 neuron279_1 (
      .a(input_layer[1212]),
      .b(input_layer[888]),
      .c(input_layer[89]),
      .d(input_layer[181]),
      .e(input_layer[100]),
      .y(Y[279]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron280_1
  function_42 neuron280_1 (
      .a(input_layer[1000]),
      .b(input_layer[476]),
      .c(input_layer[1128]),
      .d(input_layer[1112]),
      .y(Y[280]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_134 for neuron281_1
  function_134 neuron281_1 (
      .a(input_layer[1142]),
      .b(input_layer[778]),
      .c(input_layer[515]),
      .d(input_layer[757]),
      .e(input_layer[307]),
      .f(input_layer[1280]),
      .y(Y[281]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron282_1
  function_135 neuron282_1 (
      .a(~input_layer[611]),
      .b(input_layer[1470]),
      .c(~input_layer[580]),
      .d(input_layer[1236]),
      .e(input_layer[451]),
      .y(Y[282]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron283_1
  function_85 neuron283_1 (
      .a(input_layer[538]),
      .b(input_layer[566]),
      .c(input_layer[351]),
      .d(~input_layer[718]),
      .e(input_layer[1447]),
      .f(~input_layer[778]),
      .y(Y[283]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_136 for neuron284_1
  function_136 neuron284_1 (
      .a(~input_layer[1368]),
      .b(input_layer[1061]),
      .c(~input_layer[1261]),
      .d(~input_layer[1254]),
      .e(~input_layer[787]),
      .f(~input_layer[1121]),
      .y(Y[284]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron285_1
  function_78 neuron285_1 (
      .a(~input_layer[930]),
      .b(~input_layer[517]),
      .c(~input_layer[795]),
      .d(~input_layer[289]),
      .e(~input_layer[1553]),
      .f(~input_layer[335]),
      .y(Y[285]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron286_1
  function_29 neuron286_1 (
      .a(~input_layer[1250]),
      .b(~input_layer[1201]),
      .y(Y[286]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron287_1
  function_90 neuron287_1 (
      .a(input_layer[1086]),
      .b(~input_layer[373]),
      .c(~input_layer[876]),
      .d(~input_layer[1268]),
      .e(input_layer[88]),
      .y(Y[287]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron288_1
  function_11 neuron288_1 (
      .a(input_layer[577]),
      .b(~input_layer[289]),
      .c(~input_layer[1078]),
      .d(~input_layer[813]),
      .y(Y[288]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron289_1
  function_35 neuron289_1 (
      .a(~input_layer[495]),
      .b(~input_layer[498]),
      .c(~input_layer[359]),
      .d(~input_layer[98]),
      .e(~input_layer[488]),
      .y(Y[289]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_105 for neuron290_1
  function_105 neuron290_1 (
      .a(~input_layer[329]),
      .b(input_layer[365]),
      .c(input_layer[1087]),
      .d(input_layer[315]),
      .e(~input_layer[954]),
      .y(Y[290]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_137 for neuron291_1
  function_137 neuron291_1 (
      .a(~input_layer[362]),
      .b(~input_layer[1350]),
      .c(input_layer[1038]),
      .d(input_layer[219]),
      .e(input_layer[1219]),
      .y(Y[291]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron292_1
  function_106 neuron292_1 (
      .a(input_layer[792]),
      .b(~input_layer[1073]),
      .c(~input_layer[1124]),
      .d(input_layer[1329]),
      .y(Y[292]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_138 for neuron293_1
  function_138 neuron293_1 (
      .a(input_layer[440]),
      .b(~input_layer[740]),
      .c(~input_layer[1498]),
      .d(~input_layer[1369]),
      .e(~input_layer[1327]),
      .f(input_layer[1556]),
      .y(Y[293]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron294_1
  function_25 neuron294_1 (
      .a(input_layer[1030]),
      .b(~input_layer[804]),
      .c(input_layer[1050]),
      .d(input_layer[586]),
      .e(input_layer[590]),
      .y(Y[294]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron295_1
  function_42 neuron295_1 (
      .a(input_layer[1487]),
      .b(input_layer[1276]),
      .c(~input_layer[1199]),
      .d(input_layer[1296]),
      .y(Y[295]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron296_1
  function_17 neuron296_1 (
      .a(~input_layer[587]),
      .b(input_layer[1072]),
      .c(input_layer[892]),
      .y(Y[296]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron297_1
  function_29 neuron297_1 (
      .a(~input_layer[816]),
      .b(~input_layer[140]),
      .y(Y[297]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron298_1
  function_139 neuron298_1 (
      .a(input_layer[859]),
      .b(~input_layer[470]),
      .c(~input_layer[515]),
      .d(input_layer[1326]),
      .e(input_layer[633]),
      .f(~input_layer[846]),
      .y(Y[298]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_81 for neuron299_1
  function_81 neuron299_1 (
      .a(input_layer[883]),
      .b(input_layer[851]),
      .c(input_layer[850]),
      .d(input_layer[591]),
      .e(~input_layer[1543]),
      .f(input_layer[275]),
      .y(Y[299]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_140 for neuron300_1
  function_140 neuron300_1 (
      .a(~input_layer[775]),
      .b(input_layer[1246]),
      .c(~input_layer[1494]),
      .d(~input_layer[1145]),
      .e(input_layer[1163]),
      .f(~input_layer[985]),
      .y(Y[300]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron301_1
  function_119 neuron301_1 (
      .a(~input_layer[597]),
      .b(~input_layer[472]),
      .c(~input_layer[1409]),
      .d(input_layer[115]),
      .e(~input_layer[1231]),
      .y(Y[301]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_141 for neuron302_1
  function_141 neuron302_1 (
      .a(input_layer[1053]),
      .b(input_layer[695]),
      .c(input_layer[138]),
      .d(input_layer[645]),
      .e(~input_layer[569]),
      .f(~input_layer[904]),
      .y(Y[302]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron303_1
  function_16 neuron303_1 (
      .a(input_layer[597]),
      .b(~input_layer[318]),
      .y(Y[303]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron304_1
  function_26 neuron304_1 (
      .a(input_layer[637]),
      .y(Y[304]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron305_1
  function_28 neuron305_1 (
      .a(~input_layer[1418]),
      .b(~input_layer[438]),
      .c(~input_layer[931]),
      .d(~input_layer[1351]),
      .e(~input_layer[1532]),
      .f(~input_layer[1533]),
      .y(Y[305]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron306_1
  function_17 neuron306_1 (
      .a(input_layer[868]),
      .b(input_layer[1427]),
      .c(input_layer[760]),
      .y(Y[306]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron307_1
  function_60 neuron307_1 (
      .a(input_layer[1242]),
      .b(~input_layer[653]),
      .c(input_layer[298]),
      .d(input_layer[559]),
      .e(input_layer[296]),
      .y(Y[307]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_142 for neuron308_1
  function_142 neuron308_1 (
      .a(~input_layer[594]),
      .b(input_layer[632]),
      .c(~input_layer[994]),
      .d(~input_layer[233]),
      .e(~input_layer[206]),
      .f(input_layer[802]),
      .y(Y[308]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron309_1
  function_31 neuron309_1 (
      .a(~input_layer[889]),
      .b(input_layer[1117]),
      .c(~input_layer[912]),
      .d(~input_layer[859]),
      .y(Y[309]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron310_1
  function_27 neuron310_1 (
      .a(input_layer[718]),
      .b(~input_layer[274]),
      .c(~input_layer[1548]),
      .y(Y[310]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron311_1
  function_59 neuron311_1 (
      .a(~input_layer[1084]),
      .b(input_layer[232]),
      .c(input_layer[1298]),
      .d(input_layer[421]),
      .e(~input_layer[666]),
      .f(~input_layer[379]),
      .y(Y[311]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_143 for neuron312_1
  function_143 neuron312_1 (
      .a(input_layer[186]),
      .b(~input_layer[981]),
      .c(input_layer[178]),
      .d(input_layer[1393]),
      .e(input_layer[98]),
      .f(~input_layer[432]),
      .y(Y[312]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron313_1
  function_31 neuron313_1 (
      .a(input_layer[567]),
      .b(~input_layer[1311]),
      .c(input_layer[956]),
      .d(~input_layer[1114]),
      .y(Y[313]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron314_1
  function_27 neuron314_1 (
      .a(~input_layer[716]),
      .b(~input_layer[144]),
      .c(input_layer[437]),
      .y(Y[314]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron315_1
  function_100 neuron315_1 (
      .a(~input_layer[1082]),
      .b(~input_layer[795]),
      .c(~input_layer[611]),
      .d(input_layer[1155]),
      .e(input_layer[429]),
      .f(input_layer[93]),
      .y(Y[315]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron316_1
  function_27 neuron316_1 (
      .a(~input_layer[883]),
      .b(~input_layer[1475]),
      .c(input_layer[871]),
      .y(Y[316]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron317_1
  function_11 neuron317_1 (
      .a(~input_layer[943]),
      .b(~input_layer[406]),
      .c(input_layer[816]),
      .d(input_layer[85]),
      .y(Y[317]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_144 for neuron318_1
  function_144 neuron318_1 (
      .a(~input_layer[1150]),
      .b(~input_layer[1442]),
      .c(~input_layer[792]),
      .d(input_layer[1110]),
      .e(~input_layer[803]),
      .f(input_layer[1394]),
      .y(Y[318]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron319_1
  function_42 neuron319_1 (
      .a(input_layer[770]),
      .b(input_layer[803]),
      .c(input_layer[915]),
      .d(input_layer[737]),
      .y(Y[319]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron320_1
  function_42 neuron320_1 (
      .a(input_layer[972]),
      .b(input_layer[540]),
      .c(input_layer[651]),
      .d(input_layer[569]),
      .y(Y[320]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron321_1
  function_36 neuron321_1 (
      .a(input_layer[414]),
      .b(input_layer[516]),
      .c(input_layer[568]),
      .d(~input_layer[1035]),
      .e(input_layer[1531]),
      .f(input_layer[565]),
      .y(Y[321]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron322_1
  function_12 neuron322_1 (
      .a(input_layer[635]),
      .b(~input_layer[1270]),
      .c(~input_layer[907]),
      .y(Y[322]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron323_1
  function_145 neuron323_1 (
      .a(input_layer[1193]),
      .b(input_layer[571]),
      .c(~input_layer[198]),
      .d(~input_layer[827]),
      .e(~input_layer[241]),
      .y(Y[323]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron324_1
  function_55 neuron324_1 (
      .a(~input_layer[522]),
      .b(~input_layer[416]),
      .c(~input_layer[818]),
      .d(~input_layer[509]),
      .e(~input_layer[1500]),
      .y(Y[324]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron325_1
  function_120 neuron325_1 (
      .a(~input_layer[199]),
      .b(input_layer[1543]),
      .c(input_layer[551]),
      .d(input_layer[1527]),
      .e(~input_layer[883]),
      .y(Y[325]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron326_1
  function_146 neuron326_1 (
      .a(input_layer[1486]),
      .b(input_layer[846]),
      .c(~input_layer[918]),
      .d(input_layer[456]),
      .e(input_layer[915]),
      .f(input_layer[1152]),
      .y(Y[326]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron327_1
  function_26 neuron327_1 (
      .a(~input_layer[534]),
      .y(Y[327]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[328] = 1'b0;

  // instantiate function_147 for neuron329_1
  function_147 neuron329_1 (
      .a(input_layer[1390]),
      .b(~input_layer[775]),
      .c(~input_layer[1248]),
      .d(~input_layer[938]),
      .e(input_layer[666]),
      .f(~input_layer[507]),
      .y(Y[329]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron330_1
  function_148 neuron330_1 (
      .a(input_layer[624]),
      .b(~input_layer[860]),
      .c(input_layer[565]),
      .d(~input_layer[161]),
      .e(input_layer[1504]),
      .f(~input_layer[393]),
      .y(Y[330]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron331_1
  function_29 neuron331_1 (
      .a(~input_layer[415]),
      .b(~input_layer[455]),
      .y(Y[331]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron332_1
  function_74 neuron332_1 (
      .a(~input_layer[260]),
      .b(~input_layer[76]),
      .c(~input_layer[1126]),
      .d(~input_layer[1404]),
      .e(~input_layer[229]),
      .f(input_layer[1554]),
      .y(Y[332]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron333_1
  function_42 neuron333_1 (
      .a(input_layer[196]),
      .b(input_layer[643]),
      .c(input_layer[206]),
      .d(~input_layer[747]),
      .y(Y[333]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron334_1
  function_149 neuron334_1 (
      .a(input_layer[212]),
      .b(input_layer[154]),
      .c(~input_layer[1363]),
      .d(~input_layer[1167]),
      .y(Y[334]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron335_1
  function_17 neuron335_1 (
      .a(input_layer[308]),
      .b(input_layer[203]),
      .c(input_layer[1297]),
      .y(Y[335]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron336_1
  function_17 neuron336_1 (
      .a(input_layer[821]),
      .b(input_layer[1485]),
      .c(input_layer[1478]),
      .y(Y[336]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron337_1
  function_7 neuron337_1 (
      .a(input_layer[205]),
      .b(~input_layer[806]),
      .c(input_layer[513]),
      .d(~input_layer[640]),
      .y(Y[337]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_150 for neuron338_1
  function_150 neuron338_1 (
      .a(input_layer[855]),
      .b(~input_layer[1181]),
      .c(~input_layer[761]),
      .d(input_layer[666]),
      .e(input_layer[861]),
      .f(input_layer[70]),
      .y(Y[338]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron339_1
  function_3 neuron339_1 (
      .a(~input_layer[878]),
      .b(~input_layer[556]),
      .c(~input_layer[1292]),
      .d(~input_layer[367]),
      .y(Y[339]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron340_1
  function_56 neuron340_1 (
      .a(input_layer[1084]),
      .b(~input_layer[801]),
      .c(input_layer[1147]),
      .d(input_layer[716]),
      .e(input_layer[516]),
      .y(Y[340]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_151 for neuron341_1
  function_151 neuron341_1 (
      .a(~input_layer[202]),
      .b(input_layer[416]),
      .c(~input_layer[579]),
      .d(input_layer[1122]),
      .e(~input_layer[101]),
      .f(input_layer[731]),
      .y(Y[341]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron342_1
  function_152 neuron342_1 (
      .a(input_layer[981]),
      .b(~input_layer[797]),
      .c(input_layer[909]),
      .d(~input_layer[1548]),
      .e(~input_layer[131]),
      .y(Y[342]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron343_1
  function_130 neuron343_1 (
      .a(input_layer[253]),
      .b(~input_layer[739]),
      .c(input_layer[1163]),
      .d(~input_layer[794]),
      .e(input_layer[1268]),
      .f(input_layer[879]),
      .y(Y[343]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[344] = 1'b0;

  // instantiate function_24 for neuron345_1
  function_24 neuron345_1 (
      .a(input_layer[921]),
      .b(~input_layer[1045]),
      .c(~input_layer[360]),
      .y(Y[345]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_153 for neuron346_1
  function_153 neuron346_1 (
      .a(input_layer[815]),
      .b(~input_layer[947]),
      .c(input_layer[77]),
      .d(input_layer[1446]),
      .e(~input_layer[1100]),
      .f(input_layer[727]),
      .y(Y[346]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron347_1
  function_154 neuron347_1 (
      .a(~input_layer[1427]),
      .b(~input_layer[1157]),
      .c(input_layer[648]),
      .d(input_layer[266]),
      .e(input_layer[670]),
      .f(input_layer[95]),
      .y(Y[347]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron348_1
  function_3 neuron348_1 (
      .a(~input_layer[931]),
      .b(~input_layer[999]),
      .c(~input_layer[581]),
      .d(input_layer[700]),
      .y(Y[348]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron349_1
  function_155 neuron349_1 (
      .a(~input_layer[885]),
      .b(~input_layer[621]),
      .c(~input_layer[1158]),
      .d(~input_layer[663]),
      .e(~input_layer[288]),
      .f(~input_layer[731]),
      .y(Y[349]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron350_1
  function_30 neuron350_1 (
      .a(input_layer[695]),
      .b(input_layer[183]),
      .c(~input_layer[1036]),
      .d(input_layer[1374]),
      .y(Y[350]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron351_1
  function_24 neuron351_1 (
      .a(input_layer[369]),
      .b(~input_layer[210]),
      .c(input_layer[406]),
      .y(Y[351]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron352_1
  function_29 neuron352_1 (
      .a(~input_layer[1298]),
      .b(input_layer[929]),
      .y(Y[352]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron353_1
  function_29 neuron353_1 (
      .a(~input_layer[772]),
      .b(~input_layer[79]),
      .y(Y[353]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron354_1
  function_156 neuron354_1 (
      .a(~input_layer[809]),
      .b(~input_layer[1218]),
      .c(input_layer[1428]),
      .d(~input_layer[1086]),
      .e(input_layer[1334]),
      .f(input_layer[398]),
      .y(Y[354]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron355_1
  function_29 neuron355_1 (
      .a(~input_layer[636]),
      .b(~input_layer[465]),
      .y(Y[355]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron356_1
  function_42 neuron356_1 (
      .a(input_layer[666]),
      .b(input_layer[1292]),
      .c(~input_layer[584]),
      .d(input_layer[1091]),
      .y(Y[356]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron357_1
  function_157 neuron357_1 (
      .a(input_layer[923]),
      .b(~input_layer[971]),
      .c(~input_layer[288]),
      .d(~input_layer[1144]),
      .e(input_layer[1395]),
      .f(~input_layer[1251]),
      .y(Y[357]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron358_1
  function_119 neuron358_1 (
      .a(input_layer[650]),
      .b(~input_layer[676]),
      .c(~input_layer[84]),
      .d(input_layer[1413]),
      .e(~input_layer[172]),
      .y(Y[358]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_158 for neuron359_1
  function_158 neuron359_1 (
      .a(input_layer[684]),
      .b(input_layer[694]),
      .c(input_layer[510]),
      .d(~input_layer[852]),
      .e(input_layer[1237]),
      .f(~input_layer[656]),
      .y(Y[359]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron360_1
  function_39 neuron360_1 (
      .a(~input_layer[967]),
      .b(input_layer[487]),
      .c(input_layer[657]),
      .y(Y[360]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron361_1
  function_46 neuron361_1 (
      .a(input_layer[659]),
      .b(input_layer[654]),
      .c(input_layer[202]),
      .d(~input_layer[563]),
      .e(~input_layer[568]),
      .y(Y[361]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron362_1
  function_27 neuron362_1 (
      .a(~input_layer[474]),
      .b(~input_layer[1182]),
      .c(input_layer[690]),
      .y(Y[362]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron363_1
  function_25 neuron363_1 (
      .a(input_layer[147]),
      .b(input_layer[1180]),
      .c(~input_layer[574]),
      .d(input_layer[945]),
      .e(~input_layer[640]),
      .y(Y[363]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron364_1
  function_27 neuron364_1 (
      .a(~input_layer[828]),
      .b(input_layer[1108]),
      .c(~input_layer[1482]),
      .y(Y[364]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron365_1
  function_17 neuron365_1 (
      .a(input_layer[549]),
      .b(input_layer[529]),
      .c(input_layer[419]),
      .y(Y[365]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_159 for neuron366_1
  function_159 neuron366_1 (
      .a(~input_layer[422]),
      .b(input_layer[324]),
      .c(input_layer[430]),
      .d(~input_layer[834]),
      .e(~input_layer[1223]),
      .f(~input_layer[1507]),
      .y(Y[366]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[367] = 1'b0;

  // instantiate function_160 for neuron368_1
  function_160 neuron368_1 (
      .a(input_layer[662]),
      .b(~input_layer[1125]),
      .c(~input_layer[703]),
      .d(~input_layer[458]),
      .e(~input_layer[343]),
      .f(~input_layer[1046]),
      .y(Y[368]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_161 for neuron369_1
  function_161 neuron369_1 (
      .a(~input_layer[1014]),
      .b(~input_layer[1004]),
      .c(input_layer[859]),
      .d(input_layer[1548]),
      .e(~input_layer[1325]),
      .f(~input_layer[1200]),
      .y(Y[369]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron370_1
  function_149 neuron370_1 (
      .a(input_layer[882]),
      .b(~input_layer[1004]),
      .c(~input_layer[373]),
      .d(~input_layer[605]),
      .y(Y[370]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron371_1
  function_48 neuron371_1 (
      .a(input_layer[198]),
      .b(input_layer[237]),
      .c(input_layer[1384]),
      .d(~input_layer[1361]),
      .e(input_layer[559]),
      .y(Y[371]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron372_1
  function_162 neuron372_1 (
      .a(~input_layer[915]),
      .b(input_layer[648]),
      .c(input_layer[556]),
      .d(~input_layer[313]),
      .e(input_layer[402]),
      .f(input_layer[921]),
      .y(Y[372]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron373_1
  function_154 neuron373_1 (
      .a(~input_layer[1088]),
      .b(~input_layer[262]),
      .c(~input_layer[562]),
      .d(~input_layer[1338]),
      .e(input_layer[21]),
      .f(input_layer[105]),
      .y(Y[373]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron374_1
  function_7 neuron374_1 (
      .a(input_layer[552]),
      .b(~input_layer[644]),
      .c(input_layer[1146]),
      .d(~input_layer[243]),
      .y(Y[374]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron375_1
  function_26 neuron375_1 (
      .a(input_layer[810]),
      .y(Y[375]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron376_1
  function_55 neuron376_1 (
      .a(~input_layer[1539]),
      .b(~input_layer[1255]),
      .c(~input_layer[240]),
      .d(input_layer[491]),
      .e(input_layer[1387]),
      .y(Y[376]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron377_1
  function_17 neuron377_1 (
      .a(input_layer[1127]),
      .b(input_layer[1418]),
      .c(~input_layer[747]),
      .y(Y[377]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron378_1
  function_112 neuron378_1 (
      .a(input_layer[651]),
      .b(~input_layer[384]),
      .c(~input_layer[1415]),
      .d(~input_layer[850]),
      .e(input_layer[1124]),
      .f(input_layer[670]),
      .y(Y[378]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron379_1
  function_48 neuron379_1 (
      .a(~input_layer[1030]),
      .b(input_layer[857]),
      .c(input_layer[1393]),
      .d(input_layer[1339]),
      .e(input_layer[1435]),
      .y(Y[379]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_163 for neuron380_1
  function_163 neuron380_1 (
      .a(input_layer[758]),
      .b(~input_layer[967]),
      .c(~input_layer[1140]),
      .d(input_layer[233]),
      .e(input_layer[536]),
      .y(Y[380]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron381_1
  function_39 neuron381_1 (
      .a(input_layer[1266]),
      .b(~input_layer[1534]),
      .c(~input_layer[965]),
      .y(Y[381]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_164 for neuron382_1
  function_164 neuron382_1 (
      .a(~input_layer[364]),
      .b(~input_layer[892]),
      .c(input_layer[1041]),
      .d(input_layer[475]),
      .e(input_layer[57]),
      .f(input_layer[1262]),
      .y(Y[382]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron383_1
  function_123 neuron383_1 (
      .a(input_layer[196]),
      .b(~input_layer[795]),
      .c(~input_layer[342]),
      .d(input_layer[587]),
      .y(Y[383]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron384_1
  function_27 neuron384_1 (
      .a(~input_layer[405]),
      .b(~input_layer[313]),
      .c(~input_layer[1298]),
      .y(Y[384]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron385_1
  function_148 neuron385_1 (
      .a(input_layer[882]),
      .b(input_layer[1543]),
      .c(~input_layer[363]),
      .d(input_layer[230]),
      .e(input_layer[615]),
      .f(input_layer[842]),
      .y(Y[385]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron386_1
  function_6 neuron386_1 (
      .a(~input_layer[1430]),
      .b(~input_layer[1503]),
      .c(input_layer[218]),
      .d(input_layer[125]),
      .e(input_layer[338]),
      .f(input_layer[392]),
      .y(Y[386]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron387_1
  function_165 neuron387_1 (
      .a(input_layer[311]),
      .b(~input_layer[849]),
      .c(~input_layer[1429]),
      .d(input_layer[1099]),
      .e(~input_layer[1341]),
      .y(Y[387]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_166 for neuron388_1
  function_166 neuron388_1 (
      .a(~input_layer[717]),
      .b(~input_layer[1026]),
      .c(input_layer[795]),
      .d(input_layer[570]),
      .e(~input_layer[1520]),
      .f(input_layer[1400]),
      .y(Y[388]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron389_1
  function_7 neuron389_1 (
      .a(input_layer[1476]),
      .b(~input_layer[585]),
      .c(~input_layer[667]),
      .d(input_layer[446]),
      .y(Y[389]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron390_1
  function_28 neuron390_1 (
      .a(~input_layer[835]),
      .b(~input_layer[567]),
      .c(~input_layer[265]),
      .d(~input_layer[1261]),
      .e(~input_layer[732]),
      .f(~input_layer[287]),
      .y(Y[390]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron391_1
  function_27 neuron391_1 (
      .a(~input_layer[1369]),
      .b(~input_layer[1271]),
      .c(~input_layer[849]),
      .y(Y[391]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron392_1
  function_27 neuron392_1 (
      .a(~input_layer[712]),
      .b(~input_layer[236]),
      .c(input_layer[376]),
      .y(Y[392]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron393_1
  function_167 neuron393_1 (
      .a(input_layer[1056]),
      .b(input_layer[693]),
      .c(input_layer[586]),
      .d(input_layer[1479]),
      .e(~input_layer[961]),
      .y(Y[393]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron394_1
  function_29 neuron394_1 (
      .a(~input_layer[1022]),
      .b(~input_layer[1244]),
      .y(Y[394]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_168 for neuron395_1
  function_168 neuron395_1 (
      .a(~input_layer[801]),
      .b(input_layer[702]),
      .c(input_layer[361]),
      .d(~input_layer[382]),
      .e(input_layer[547]),
      .f(input_layer[1005]),
      .y(Y[395]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron396_1
  function_169 neuron396_1 (
      .a(~input_layer[1428]),
      .b(~input_layer[488]),
      .c(input_layer[155]),
      .d(input_layer[915]),
      .e(input_layer[930]),
      .f(input_layer[1454]),
      .y(Y[396]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron397_1
  function_170 neuron397_1 (
      .a(~input_layer[1481]),
      .b(input_layer[1374]),
      .c(~input_layer[160]),
      .d(input_layer[439]),
      .e(input_layer[1078]),
      .f(input_layer[1204]),
      .y(Y[397]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron398_1
  function_87 neuron398_1 (
      .a(input_layer[299]),
      .b(~input_layer[718]),
      .c(input_layer[1098]),
      .d(input_layer[895]),
      .e(~input_layer[395]),
      .y(Y[398]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron399_1
  function_0 neuron399_1 (
      .a(~input_layer[492]),
      .b(~input_layer[372]),
      .c(~input_layer[267]),
      .d(~input_layer[209]),
      .e(~input_layer[139]),
      .y(Y[399]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron400_1
  function_48 neuron400_1 (
      .a(input_layer[556]),
      .b(input_layer[1081]),
      .c(input_layer[1221]),
      .d(input_layer[780]),
      .e(~input_layer[1377]),
      .y(Y[400]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron401_1
  function_106 neuron401_1 (
      .a(input_layer[370]),
      .b(input_layer[515]),
      .c(input_layer[468]),
      .d(~input_layer[976]),
      .y(Y[401]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron402_1
  function_7 neuron402_1 (
      .a(~input_layer[694]),
      .b(input_layer[734]),
      .c(input_layer[1420]),
      .d(~input_layer[1096]),
      .y(Y[402]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron403_1
  function_78 neuron403_1 (
      .a(~input_layer[664]),
      .b(~input_layer[241]),
      .c(~input_layer[1243]),
      .d(~input_layer[154]),
      .e(input_layer[395]),
      .f(input_layer[486]),
      .y(Y[403]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_171 for neuron404_1
  function_171 neuron404_1 (
      .a(input_layer[1184]),
      .b(~input_layer[743]),
      .c(~input_layer[1534]),
      .d(input_layer[570]),
      .e(~input_layer[142]),
      .f(input_layer[1380]),
      .y(Y[404]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron405_1
  function_87 neuron405_1 (
      .a(input_layer[1432]),
      .b(~input_layer[1083]),
      .c(input_layer[955]),
      .d(~input_layer[895]),
      .e(input_layer[410]),
      .y(Y[405]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron406_1
  function_19 neuron406_1 (
      .a(~input_layer[207]),
      .b(~input_layer[868]),
      .c(~input_layer[191]),
      .d(input_layer[564]),
      .y(Y[406]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron407_1
  function_59 neuron407_1 (
      .a(input_layer[1030]),
      .b(~input_layer[590]),
      .c(input_layer[1170]),
      .d(input_layer[1034]),
      .e(~input_layer[1250]),
      .f(~input_layer[1154]),
      .y(Y[407]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron408_1
  function_26 neuron408_1 (
      .a(~input_layer[762]),
      .y(Y[408]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron409_1
  function_172 neuron409_1 (
      .a(~input_layer[1313]),
      .b(~input_layer[455]),
      .c(input_layer[76]),
      .d(~input_layer[1465]),
      .e(~input_layer[451]),
      .f(~input_layer[450]),
      .y(Y[409]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron410_1
  function_24 neuron410_1 (
      .a(~input_layer[642]),
      .b(input_layer[197]),
      .c(~input_layer[1532]),
      .y(Y[410]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron411_1
  function_27 neuron411_1 (
      .a(~input_layer[1071]),
      .b(~input_layer[983]),
      .c(~input_layer[622]),
      .y(Y[411]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron412_1
  function_27 neuron412_1 (
      .a(~input_layer[420]),
      .b(~input_layer[1484]),
      .c(~input_layer[1055]),
      .y(Y[412]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[413] = 1'b1;

  // instantiate function_26 for neuron414_1
  function_26 neuron414_1 (
      .a(~input_layer[867]),
      .y(Y[414]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron415_1
  function_84 neuron415_1 (
      .a(~input_layer[965]),
      .b(~input_layer[711]),
      .c(input_layer[1247]),
      .d(~input_layer[1250]),
      .e(~input_layer[256]),
      .y(Y[415]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_173 for neuron416_1
  function_173 neuron416_1 (
      .a(~input_layer[1028]),
      .b(input_layer[1305]),
      .c(~input_layer[1003]),
      .d(~input_layer[804]),
      .e(~input_layer[85]),
      .y(Y[416]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron417_1
  function_42 neuron417_1 (
      .a(input_layer[349]),
      .b(input_layer[887]),
      .c(input_layer[942]),
      .d(input_layer[1257]),
      .y(Y[417]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron418_1
  function_3 neuron418_1 (
      .a(~input_layer[359]),
      .b(~input_layer[516]),
      .c(~input_layer[779]),
      .d(~input_layer[1306]),
      .y(Y[418]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron419_1
  function_47 neuron419_1 (
      .a(input_layer[1220]),
      .b(input_layer[197]),
      .c(input_layer[1103]),
      .d(input_layer[127]),
      .e(input_layer[983]),
      .y(Y[419]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron420_1
  function_26 neuron420_1 (
      .a(input_layer[144]),
      .y(Y[420]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron421_1
  function_36 neuron421_1 (
      .a(input_layer[1053]),
      .b(input_layer[186]),
      .c(input_layer[834]),
      .d(input_layer[1012]),
      .e(input_layer[1280]),
      .f(input_layer[1285]),
      .y(Y[421]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron422_1
  function_24 neuron422_1 (
      .a(input_layer[546]),
      .b(~input_layer[128]),
      .c(~input_layer[1045]),
      .y(Y[422]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron423_1
  function_67 neuron423_1 (
      .a(~input_layer[579]),
      .b(~input_layer[772]),
      .c(~input_layer[1482]),
      .d(~input_layer[420]),
      .e(~input_layer[1537]),
      .y(Y[423]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron424_1
  function_3 neuron424_1 (
      .a(~input_layer[524]),
      .b(~input_layer[1126]),
      .c(~input_layer[929]),
      .d(~input_layer[1295]),
      .y(Y[424]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron425_1
  function_26 neuron425_1 (
      .a(input_layer[1202]),
      .y(Y[425]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron426_1
  function_31 neuron426_1 (
      .a(input_layer[948]),
      .b(~input_layer[654]),
      .c(~input_layer[849]),
      .d(~input_layer[1215]),
      .y(Y[426]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_174 for neuron427_1
  function_174 neuron427_1 (
      .a(~input_layer[1137]),
      .b(input_layer[211]),
      .c(input_layer[877]),
      .d(~input_layer[241]),
      .e(input_layer[751]),
      .f(input_layer[288]),
      .y(Y[427]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron428_1
  function_175 neuron428_1 (
      .a(input_layer[444]),
      .b(input_layer[419]),
      .c(input_layer[1261]),
      .d(~input_layer[1553]),
      .e(~input_layer[999]),
      .f(input_layer[1503]),
      .y(Y[428]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron429_1
  function_19 neuron429_1 (
      .a(~input_layer[384]),
      .b(~input_layer[699]),
      .c(input_layer[1370]),
      .d(~input_layer[900]),
      .y(Y[429]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron430_1
  function_55 neuron430_1 (
      .a(~input_layer[150]),
      .b(~input_layer[1158]),
      .c(~input_layer[256]),
      .d(~input_layer[1124]),
      .e(input_layer[552]),
      .y(Y[430]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron431_1
  function_24 neuron431_1 (
      .a(~input_layer[740]),
      .b(input_layer[930]),
      .c(~input_layer[491]),
      .y(Y[431]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron432_1
  function_17 neuron432_1 (
      .a(~input_layer[1022]),
      .b(input_layer[212]),
      .c(input_layer[1546]),
      .y(Y[432]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_164 for neuron433_1
  function_164 neuron433_1 (
      .a(~input_layer[591]),
      .b(~input_layer[1187]),
      .c(input_layer[601]),
      .d(input_layer[1539]),
      .e(~input_layer[1045]),
      .f(~input_layer[1178]),
      .y(Y[433]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron434_1
  function_1 neuron434_1 (
      .a(~input_layer[925]),
      .b(input_layer[643]),
      .c(~input_layer[1528]),
      .d(~input_layer[961]),
      .y(Y[434]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron435_1
  function_27 neuron435_1 (
      .a(~input_layer[382]),
      .b(input_layer[1090]),
      .c(~input_layer[907]),
      .y(Y[435]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron436_1
  function_42 neuron436_1 (
      .a(input_layer[1226]),
      .b(input_layer[665]),
      .c(~input_layer[804]),
      .d(input_layer[481]),
      .y(Y[436]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_176 for neuron437_1
  function_176 neuron437_1 (
      .a(input_layer[1181]),
      .b(input_layer[455]),
      .c(~input_layer[970]),
      .d(~input_layer[1040]),
      .e(~input_layer[822]),
      .f(input_layer[231]),
      .y(Y[437]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_102 for neuron438_1
  function_102 neuron438_1 (
      .a(~input_layer[862]),
      .b(~input_layer[310]),
      .c(input_layer[710]),
      .d(~input_layer[1013]),
      .e(~input_layer[1266]),
      .f(input_layer[487]),
      .y(Y[438]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron439_1
  function_123 neuron439_1 (
      .a(input_layer[602]),
      .b(input_layer[258]),
      .c(input_layer[431]),
      .d(~input_layer[435]),
      .y(Y[439]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron440_1
  function_29 neuron440_1 (
      .a(~input_layer[641]),
      .b(~input_layer[1261]),
      .y(Y[440]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron441_1
  function_16 neuron441_1 (
      .a(input_layer[272]),
      .b(~input_layer[1333]),
      .y(Y[441]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron442_1
  function_74 neuron442_1 (
      .a(~input_layer[879]),
      .b(input_layer[471]),
      .c(~input_layer[847]),
      .d(~input_layer[646]),
      .e(~input_layer[817]),
      .f(~input_layer[119]),
      .y(Y[442]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron443_1
  function_63 neuron443_1 (
      .a(~input_layer[1300]),
      .b(input_layer[147]),
      .c(input_layer[886]),
      .d(~input_layer[666]),
      .e(input_layer[181]),
      .y(Y[443]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_177 for neuron444_1
  function_177 neuron444_1 (
      .a(~input_layer[139]),
      .b(input_layer[766]),
      .c(input_layer[652]),
      .d(input_layer[1369]),
      .e(input_layer[1525]),
      .y(Y[444]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron445_1
  function_167 neuron445_1 (
      .a(input_layer[209]),
      .b(input_layer[1388]),
      .c(~input_layer[398]),
      .d(input_layer[503]),
      .e(~input_layer[1522]),
      .y(Y[445]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_178 for neuron446_1
  function_178 neuron446_1 (
      .a(~input_layer[1034]),
      .b(input_layer[360]),
      .c(~input_layer[1472]),
      .d(~input_layer[86]),
      .e(input_layer[647]),
      .f(input_layer[1005]),
      .y(Y[446]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron447_1
  function_42 neuron447_1 (
      .a(input_layer[1423]),
      .b(input_layer[496]),
      .c(input_layer[963]),
      .d(input_layer[653]),
      .y(Y[447]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron448_1
  function_12 neuron448_1 (
      .a(input_layer[577]),
      .b(~input_layer[308]),
      .c(~input_layer[1299]),
      .y(Y[448]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron449_1
  function_8 neuron449_1 (
      .a(input_layer[478]),
      .b(input_layer[1492]),
      .c(~input_layer[692]),
      .d(input_layer[1079]),
      .y(Y[449]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron450_1
  function_179 neuron450_1 (
      .a(~input_layer[697]),
      .b(~input_layer[554]),
      .c(~input_layer[775]),
      .d(input_layer[931]),
      .e(input_layer[1533]),
      .y(Y[450]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_180 for neuron451_1
  function_180 neuron451_1 (
      .a(input_layer[867]),
      .b(~input_layer[306]),
      .c(input_layer[568]),
      .d(~input_layer[1077]),
      .e(~input_layer[1132]),
      .f(~input_layer[1219]),
      .y(Y[451]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron452_1
  function_12 neuron452_1 (
      .a(input_layer[699]),
      .b(input_layer[734]),
      .c(~input_layer[471]),
      .y(Y[452]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron453_1
  function_181 neuron453_1 (
      .a(input_layer[305]),
      .b(input_layer[832]),
      .c(~input_layer[1433]),
      .d(input_layer[1470]),
      .e(~input_layer[881]),
      .y(Y[453]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_182 for neuron454_1
  function_182 neuron454_1 (
      .a(input_layer[521]),
      .b(~input_layer[990]),
      .c(~input_layer[256]),
      .d(~input_layer[1197]),
      .e(~input_layer[850]),
      .f(~input_layer[1072]),
      .y(Y[454]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron455_1
  function_31 neuron455_1 (
      .a(input_layer[441]),
      .b(~input_layer[905]),
      .c(input_layer[607]),
      .d(~input_layer[890]),
      .y(Y[455]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron456_1
  function_183 neuron456_1 (
      .a(~input_layer[863]),
      .b(input_layer[542]),
      .c(input_layer[1282]),
      .d(~input_layer[243]),
      .e(input_layer[1063]),
      .f(input_layer[1062]),
      .y(Y[456]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron457_1
  function_46 neuron457_1 (
      .a(input_layer[973]),
      .b(input_layer[213]),
      .c(input_layer[1112]),
      .d(~input_layer[252]),
      .e(input_layer[179]),
      .y(Y[457]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron458_1
  function_92 neuron458_1 (
      .a(input_layer[1269]),
      .b(input_layer[664]),
      .c(input_layer[1027]),
      .d(~input_layer[933]),
      .e(~input_layer[816]),
      .f(input_layer[1096]),
      .y(Y[458]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_184 for neuron459_1
  function_184 neuron459_1 (
      .a(input_layer[1183]),
      .b(~input_layer[1083]),
      .c(~input_layer[131]),
      .d(~input_layer[83]),
      .e(input_layer[1262]),
      .y(Y[459]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_185 for neuron460_1
  function_185 neuron460_1 (
      .a(input_layer[977]),
      .b(~input_layer[1267]),
      .c(input_layer[814]),
      .d(input_layer[209]),
      .e(~input_layer[939]),
      .f(input_layer[200]),
      .y(Y[460]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron461_1
  function_25 neuron461_1 (
      .a(input_layer[1437]),
      .b(input_layer[491]),
      .c(input_layer[370]),
      .d(input_layer[1322]),
      .e(input_layer[1217]),
      .y(Y[461]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron462_1
  function_186 neuron462_1 (
      .a(~input_layer[721]),
      .b(input_layer[386]),
      .c(input_layer[1164]),
      .d(~input_layer[642]),
      .y(Y[462]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron463_1
  function_19 neuron463_1 (
      .a(~input_layer[1108]),
      .b(~input_layer[1135]),
      .c(input_layer[882]),
      .d(~input_layer[179]),
      .y(Y[463]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron464_1
  function_67 neuron464_1 (
      .a(~input_layer[1481]),
      .b(~input_layer[947]),
      .c(~input_layer[1422]),
      .d(~input_layer[483]),
      .e(~input_layer[1143]),
      .y(Y[464]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron465_1
  function_16 neuron465_1 (
      .a(input_layer[1247]),
      .b(~input_layer[857]),
      .y(Y[465]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron466_1
  function_67 neuron466_1 (
      .a(~input_layer[1252]),
      .b(~input_layer[1075]),
      .c(~input_layer[89]),
      .d(~input_layer[1222]),
      .e(~input_layer[205]),
      .y(Y[466]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron467_1
  function_106 neuron467_1 (
      .a(input_layer[438]),
      .b(input_layer[1435]),
      .c(~input_layer[1129]),
      .d(~input_layer[1189]),
      .y(Y[467]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron468_1
  function_47 neuron468_1 (
      .a(input_layer[932]),
      .b(input_layer[966]),
      .c(input_layer[941]),
      .d(input_layer[1227]),
      .e(input_layer[156]),
      .y(Y[468]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_187 for neuron469_1
  function_187 neuron469_1 (
      .a(input_layer[510]),
      .b(input_layer[537]),
      .c(~input_layer[1269]),
      .d(~input_layer[1004]),
      .e(~input_layer[689]),
      .f(~input_layer[726]),
      .y(Y[469]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron470_1
  function_188 neuron470_1 (
      .a(~input_layer[578]),
      .b(input_layer[452]),
      .c(~input_layer[1224]),
      .d(~input_layer[1482]),
      .e(~input_layer[1228]),
      .f(~input_layer[1172]),
      .y(Y[470]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron471_1
  function_128 neuron471_1 (
      .a(~input_layer[430]),
      .b(input_layer[146]),
      .c(input_layer[944]),
      .d(~input_layer[1351]),
      .y(Y[471]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron472_1
  function_84 neuron472_1 (
      .a(input_layer[1372]),
      .b(~input_layer[1294]),
      .c(~input_layer[219]),
      .d(~input_layer[512]),
      .e(~input_layer[1462]),
      .y(Y[472]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron473_1
  function_3 neuron473_1 (
      .a(~input_layer[495]),
      .b(~input_layer[1261]),
      .c(~input_layer[396]),
      .d(~input_layer[1280]),
      .y(Y[473]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron474_1
  function_146 neuron474_1 (
      .a(input_layer[577]),
      .b(input_layer[1259]),
      .c(~input_layer[916]),
      .d(~input_layer[1092]),
      .e(input_layer[679]),
      .f(input_layer[616]),
      .y(Y[474]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron475_1
  function_36 neuron475_1 (
      .a(input_layer[658]),
      .b(input_layer[1154]),
      .c(input_layer[241]),
      .d(input_layer[399]),
      .e(input_layer[1408]),
      .f(input_layer[178]),
      .y(Y[475]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron476_1
  function_3 neuron476_1 (
      .a(~input_layer[1434]),
      .b(~input_layer[635]),
      .c(~input_layer[291]),
      .d(~input_layer[492]),
      .y(Y[476]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron477_1
  function_3 neuron477_1 (
      .a(~input_layer[1295]),
      .b(~input_layer[887]),
      .c(~input_layer[963]),
      .d(input_layer[663]),
      .y(Y[477]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron478_1
  function_24 neuron478_1 (
      .a(~input_layer[460]),
      .b(~input_layer[648]),
      .c(input_layer[602]),
      .y(Y[478]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_189 for neuron479_1
  function_189 neuron479_1 (
      .a(~input_layer[1192]),
      .b(~input_layer[421]),
      .c(input_layer[976]),
      .d(input_layer[637]),
      .e(~input_layer[415]),
      .f(~input_layer[372]),
      .y(Y[479]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron480_1
  function_42 neuron480_1 (
      .a(input_layer[1489]),
      .b(input_layer[991]),
      .c(input_layer[993]),
      .d(input_layer[990]),
      .y(Y[480]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_190 for neuron481_1
  function_190 neuron481_1 (
      .a(input_layer[949]),
      .b(~input_layer[701]),
      .c(input_layer[1282]),
      .d(~input_layer[567]),
      .e(~input_layer[1261]),
      .f(~input_layer[1460]),
      .y(Y[481]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron482_1
  function_0 neuron482_1 (
      .a(~input_layer[1132]),
      .b(~input_layer[1253]),
      .c(~input_layer[515]),
      .d(~input_layer[516]),
      .e(input_layer[778]),
      .y(Y[482]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_191 for neuron483_1
  function_191 neuron483_1 (
      .a(input_layer[582]),
      .b(~input_layer[234]),
      .c(~input_layer[1301]),
      .d(~input_layer[1545]),
      .e(~input_layer[452]),
      .f(~input_layer[1373]),
      .y(Y[483]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron484_1
  function_167 neuron484_1 (
      .a(input_layer[1128]),
      .b(input_layer[1386]),
      .c(~input_layer[883]),
      .d(input_layer[518]),
      .e(input_layer[1216]),
      .y(Y[484]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron485_1
  function_95 neuron485_1 (
      .a(input_layer[819]),
      .b(input_layer[1440]),
      .c(~input_layer[378]),
      .d(~input_layer[1062]),
      .y(Y[485]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron486_1
  function_26 neuron486_1 (
      .a(input_layer[483]),
      .y(Y[486]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron487_1
  function_120 neuron487_1 (
      .a(input_layer[443]),
      .b(~input_layer[535]),
      .c(input_layer[1215]),
      .d(input_layer[857]),
      .e(~input_layer[1117]),
      .y(Y[487]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron488_1
  function_192 neuron488_1 (
      .a(input_layer[490]),
      .b(~input_layer[145]),
      .c(input_layer[652]),
      .d(input_layer[1416]),
      .e(input_layer[455]),
      .f(~input_layer[657]),
      .y(Y[488]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron489_1
  function_146 neuron489_1 (
      .a(~input_layer[209]),
      .b(input_layer[377]),
      .c(input_layer[789]),
      .d(input_layer[1382]),
      .e(input_layer[1118]),
      .f(~input_layer[1140]),
      .y(Y[489]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron490_1
  function_35 neuron490_1 (
      .a(~input_layer[1244]),
      .b(input_layer[764]),
      .c(~input_layer[302]),
      .d(~input_layer[963]),
      .e(~input_layer[69]),
      .y(Y[490]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron491_1
  function_193 neuron491_1 (
      .a(input_layer[1417]),
      .b(~input_layer[303]),
      .c(input_layer[155]),
      .d(input_layer[796]),
      .e(~input_layer[778]),
      .y(Y[491]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_194 for neuron492_1
  function_194 neuron492_1 (
      .a(~input_layer[308]),
      .b(~input_layer[1551]),
      .c(input_layer[765]),
      .d(~input_layer[120]),
      .e(~input_layer[462]),
      .f(input_layer[493]),
      .y(Y[492]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron493_1
  function_0 neuron493_1 (
      .a(~input_layer[136]),
      .b(~input_layer[194]),
      .c(~input_layer[1244]),
      .d(input_layer[851]),
      .e(~input_layer[451]),
      .y(Y[493]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron494_1
  function_1 neuron494_1 (
      .a(~input_layer[1418]),
      .b(input_layer[256]),
      .c(~input_layer[649]),
      .d(~input_layer[756]),
      .y(Y[494]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron495_1
  function_97 neuron495_1 (
      .a(~input_layer[595]),
      .b(~input_layer[1275]),
      .c(input_layer[1044]),
      .d(~input_layer[1130]),
      .e(input_layer[1350]),
      .y(Y[495]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron496_1
  function_16 neuron496_1 (
      .a(input_layer[610]),
      .b(input_layer[1051]),
      .y(Y[496]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron497_1
  function_19 neuron497_1 (
      .a(~input_layer[1033]),
      .b(~input_layer[215]),
      .c(input_layer[1262]),
      .d(input_layer[960]),
      .y(Y[497]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron498_1
  function_27 neuron498_1 (
      .a(~input_layer[1113]),
      .b(~input_layer[1198]),
      .c(~input_layer[359]),
      .y(Y[498]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron499_1
  function_26 neuron499_1 (
      .a(~input_layer[1028]),
      .y(Y[499]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron500_1
  function_195 neuron500_1 (
      .a(~input_layer[692]),
      .b(input_layer[1218]),
      .c(~input_layer[794]),
      .d(input_layer[487]),
      .e(input_layer[521]),
      .y(Y[500]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron501_1
  function_172 neuron501_1 (
      .a(input_layer[1018]),
      .b(~input_layer[1530]),
      .c(~input_layer[1247]),
      .d(~input_layer[677]),
      .e(~input_layer[456]),
      .f(~input_layer[1410]),
      .y(Y[501]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron502_1
  function_186 neuron502_1 (
      .a(input_layer[757]),
      .b(~input_layer[634]),
      .c(input_layer[479]),
      .d(~input_layer[524]),
      .y(Y[502]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron503_1
  function_39 neuron503_1 (
      .a(input_layer[1129]),
      .b(~input_layer[1089]),
      .c(~input_layer[523]),
      .y(Y[503]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron504_1
  function_19 neuron504_1 (
      .a(~input_layer[772]),
      .b(~input_layer[261]),
      .c(~input_layer[749]),
      .d(input_layer[245]),
      .y(Y[504]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron505_1
  function_26 neuron505_1 (
      .a(~input_layer[692]),
      .y(Y[505]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_129 for neuron506_1
  function_129 neuron506_1 (
      .a(input_layer[741]),
      .b(~input_layer[1053]),
      .c(input_layer[802]),
      .d(input_layer[651]),
      .e(~input_layer[841]),
      .f(~input_layer[828]),
      .y(Y[506]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron507_1
  function_46 neuron507_1 (
      .a(input_layer[1362]),
      .b(input_layer[1354]),
      .c(input_layer[613]),
      .d(~input_layer[692]),
      .e(~input_layer[80]),
      .y(Y[507]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron508_1
  function_27 neuron508_1 (
      .a(~input_layer[549]),
      .b(~input_layer[994]),
      .c(~input_layer[1108]),
      .y(Y[508]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron509_1
  function_26 neuron509_1 (
      .a(input_layer[425]),
      .y(Y[509]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron510_1
  function_13 neuron510_1 (
      .a(input_layer[749]),
      .b(~input_layer[1295]),
      .c(input_layer[800]),
      .d(~input_layer[1364]),
      .y(Y[510]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_196 for neuron511_1
  function_196 neuron511_1 (
      .a(~input_layer[403]),
      .b(input_layer[915]),
      .c(input_layer[690]),
      .d(~input_layer[511]),
      .e(~input_layer[1101]),
      .f(~input_layer[1192]),
      .y(Y[511]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_197 for neuron512_1
  function_197 neuron512_1 (
      .a(input_layer[1068]),
      .b(~input_layer[916]),
      .c(~input_layer[662]),
      .d(~input_layer[1497]),
      .e(~input_layer[520]),
      .f(input_layer[503]),
      .y(Y[512]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron513_1
  function_46 neuron513_1 (
      .a(input_layer[1022]),
      .b(input_layer[971]),
      .c(~input_layer[1360]),
      .d(input_layer[552]),
      .e(input_layer[1246]),
      .y(Y[513]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_83 for neuron514_1
  function_83 neuron514_1 (
      .a(input_layer[414]),
      .b(~input_layer[154]),
      .c(input_layer[380]),
      .d(~input_layer[267]),
      .e(input_layer[309]),
      .y(Y[514]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_198 for neuron515_1
  function_198 neuron515_1 (
      .a(~input_layer[701]),
      .b(input_layer[438]),
      .c(~input_layer[1252]),
      .d(~input_layer[236]),
      .e(input_layer[456]),
      .f(~input_layer[1378]),
      .y(Y[515]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron516_1
  function_39 neuron516_1 (
      .a(input_layer[510]),
      .b(~input_layer[1325]),
      .c(input_layer[521]),
      .y(Y[516]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron517_1
  function_186 neuron517_1 (
      .a(input_layer[1543]),
      .b(input_layer[874]),
      .c(~input_layer[362]),
      .d(~input_layer[1268]),
      .y(Y[517]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron518_1
  function_193 neuron518_1 (
      .a(~input_layer[580]),
      .b(input_layer[244]),
      .c(input_layer[419]),
      .d(~input_layer[872]),
      .e(~input_layer[710]),
      .y(Y[518]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron519_1
  function_0 neuron519_1 (
      .a(~input_layer[853]),
      .b(~input_layer[905]),
      .c(~input_layer[410]),
      .d(input_layer[755]),
      .e(~input_layer[1500]),
      .y(Y[519]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron520_1
  function_195 neuron520_1 (
      .a(~input_layer[353]),
      .b(input_layer[1440]),
      .c(input_layer[127]),
      .d(input_layer[391]),
      .e(input_layer[731]),
      .y(Y[520]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron521_1
  function_31 neuron521_1 (
      .a(~input_layer[580]),
      .b(input_layer[359]),
      .c(input_layer[152]),
      .d(input_layer[1189]),
      .y(Y[521]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron522_1
  function_17 neuron522_1 (
      .a(input_layer[915]),
      .b(~input_layer[1314]),
      .c(input_layer[129]),
      .y(Y[522]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron523_1
  function_97 neuron523_1 (
      .a(~input_layer[885]),
      .b(input_layer[1328]),
      .c(~input_layer[666]),
      .d(~input_layer[591]),
      .e(input_layer[198]),
      .y(Y[523]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron524_1
  function_106 neuron524_1 (
      .a(input_layer[1326]),
      .b(input_layer[376]),
      .c(~input_layer[710]),
      .d(~input_layer[1483]),
      .y(Y[524]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_199 for neuron525_1
  function_199 neuron525_1 (
      .a(~input_layer[1386]),
      .b(~input_layer[192]),
      .c(~input_layer[1391]),
      .d(input_layer[642]),
      .e(~input_layer[1264]),
      .f(~input_layer[1522]),
      .y(Y[525]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron526_1
  function_3 neuron526_1 (
      .a(~input_layer[815]),
      .b(~input_layer[622]),
      .c(~input_layer[288]),
      .d(~input_layer[984]),
      .y(Y[526]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron527_1
  function_104 neuron527_1 (
      .a(input_layer[916]),
      .b(~input_layer[1533]),
      .c(input_layer[1282]),
      .d(~input_layer[1130]),
      .e(input_layer[1231]),
      .f(input_layer[111]),
      .y(Y[527]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron528_1
  function_96 neuron528_1 (
      .a(input_layer[1087]),
      .b(~input_layer[610]),
      .c(input_layer[827]),
      .d(input_layer[120]),
      .y(Y[528]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron529_1
  function_95 neuron529_1 (
      .a(~input_layer[940]),
      .b(input_layer[1384]),
      .c(input_layer[596]),
      .d(input_layer[354]),
      .y(Y[529]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron530_1
  function_17 neuron530_1 (
      .a(input_layer[363]),
      .b(~input_layer[1370]),
      .c(input_layer[1207]),
      .y(Y[530]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_200 for neuron531_1
  function_200 neuron531_1 (
      .a(input_layer[692]),
      .b(~input_layer[539]),
      .c(~input_layer[357]),
      .d(~input_layer[249]),
      .e(~input_layer[726]),
      .f(~input_layer[1559]),
      .y(Y[531]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron532_1
  function_1 neuron532_1 (
      .a(~input_layer[1318]),
      .b(~input_layer[142]),
      .c(input_layer[892]),
      .d(input_layer[302]),
      .y(Y[532]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron533_1
  function_89 neuron533_1 (
      .a(input_layer[1190]),
      .b(~input_layer[983]),
      .c(~input_layer[980]),
      .d(~input_layer[792]),
      .e(input_layer[671]),
      .y(Y[533]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron534_1
  function_167 neuron534_1 (
      .a(input_layer[1481]),
      .b(input_layer[292]),
      .c(input_layer[1466]),
      .d(~input_layer[1022]),
      .e(~input_layer[596]),
      .y(Y[534]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron535_1
  function_12 neuron535_1 (
      .a(input_layer[639]),
      .b(~input_layer[366]),
      .c(~input_layer[985]),
      .y(Y[535]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron536_1
  function_17 neuron536_1 (
      .a(input_layer[515]),
      .b(input_layer[1369]),
      .c(~input_layer[700]),
      .y(Y[536]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron537_1
  function_3 neuron537_1 (
      .a(~input_layer[1381]),
      .b(~input_layer[545]),
      .c(~input_layer[550]),
      .d(~input_layer[1182]),
      .y(Y[537]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron538_1
  function_12 neuron538_1 (
      .a(input_layer[940]),
      .b(~input_layer[534]),
      .c(input_layer[249]),
      .y(Y[538]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron539_1
  function_0 neuron539_1 (
      .a(~input_layer[251]),
      .b(~input_layer[296]),
      .c(~input_layer[293]),
      .d(input_layer[1390]),
      .e(~input_layer[992]),
      .y(Y[539]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron540_1
  function_47 neuron540_1 (
      .a(input_layer[1090]),
      .b(~input_layer[1012]),
      .c(input_layer[1355]),
      .d(~input_layer[1407]),
      .e(~input_layer[1063]),
      .y(Y[540]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron541_1
  function_18 neuron541_1 (
      .a(input_layer[237]),
      .b(~input_layer[1135]),
      .c(~input_layer[434]),
      .d(~input_layer[1311]),
      .e(~input_layer[447]),
      .y(Y[541]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron542_1
  function_17 neuron542_1 (
      .a(~input_layer[703]),
      .b(input_layer[1435]),
      .c(input_layer[859]),
      .y(Y[542]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_201 for neuron543_1
  function_201 neuron543_1 (
      .a(input_layer[709]),
      .b(~input_layer[375]),
      .c(~input_layer[833]),
      .d(~input_layer[427]),
      .e(~input_layer[1211]),
      .f(~input_layer[895]),
      .y(Y[543]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron544_1
  function_42 neuron544_1 (
      .a(input_layer[1368]),
      .b(input_layer[606]),
      .c(~input_layer[972]),
      .d(~input_layer[1024]),
      .y(Y[544]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron545_1
  function_90 neuron545_1 (
      .a(~input_layer[328]),
      .b(~input_layer[1086]),
      .c(~input_layer[773]),
      .d(input_layer[1389]),
      .e(input_layer[1415]),
      .y(Y[545]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron546_1
  function_120 neuron546_1 (
      .a(input_layer[608]),
      .b(~input_layer[905]),
      .c(input_layer[143]),
      .d(~input_layer[771]),
      .e(input_layer[1501]),
      .y(Y[546]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron547_1
  function_202 neuron547_1 (
      .a(~input_layer[441]),
      .b(~input_layer[1365]),
      .c(input_layer[301]),
      .d(~input_layer[147]),
      .e(~input_layer[1389]),
      .f(input_layer[1228]),
      .y(Y[547]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron548_1
  function_54 neuron548_1 (
      .a(input_layer[1317]),
      .b(input_layer[1388]),
      .c(~input_layer[239]),
      .d(input_layer[503]),
      .e(~input_layer[453]),
      .f(~input_layer[765]),
      .y(Y[548]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron549_1
  function_91 neuron549_1 (
      .a(~input_layer[888]),
      .b(~input_layer[824]),
      .c(input_layer[1171]),
      .d(input_layer[455]),
      .e(input_layer[554]),
      .y(Y[549]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_203 for neuron550_1
  function_203 neuron550_1 (
      .a(input_layer[1075]),
      .b(input_layer[292]),
      .c(~input_layer[735]),
      .d(~input_layer[90]),
      .e(~input_layer[789]),
      .f(input_layer[340]),
      .y(Y[550]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_204 for neuron551_1
  function_204 neuron551_1 (
      .a(input_layer[137]),
      .b(~input_layer[1184]),
      .c(input_layer[477]),
      .d(~input_layer[1171]),
      .e(~input_layer[598]),
      .f(~input_layer[356]),
      .y(Y[551]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron552_1
  function_132 neuron552_1 (
      .a(input_layer[459]),
      .b(input_layer[243]),
      .c(input_layer[1533]),
      .d(~input_layer[741]),
      .e(~input_layer[315]),
      .f(~input_layer[33]),
      .y(Y[552]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_205 for neuron553_1
  function_205 neuron553_1 (
      .a(~input_layer[1474]),
      .b(~input_layer[1388]),
      .c(input_layer[459]),
      .d(~input_layer[471]),
      .e(input_layer[1149]),
      .f(input_layer[1341]),
      .y(Y[553]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron554_1
  function_154 neuron554_1 (
      .a(~input_layer[1219]),
      .b(~input_layer[192]),
      .c(~input_layer[191]),
      .d(input_layer[432]),
      .e(input_layer[430]),
      .f(input_layer[1066]),
      .y(Y[554]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_206 for neuron555_1
  function_206 neuron555_1 (
      .a(~input_layer[1322]),
      .b(~input_layer[1328]),
      .c(input_layer[994]),
      .d(input_layer[700]),
      .e(input_layer[27]),
      .f(input_layer[220]),
      .y(Y[555]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_207 for neuron556_1
  function_207 neuron556_1 (
      .a(input_layer[1028]),
      .b(~input_layer[400]),
      .c(input_layer[890]),
      .d(input_layer[1393]),
      .e(~input_layer[1101]),
      .f(input_layer[875]),
      .y(Y[556]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_208 for neuron557_1
  function_208 neuron557_1 (
      .a(input_layer[295]),
      .b(input_layer[513]),
      .c(input_layer[243]),
      .d(~input_layer[886]),
      .e(input_layer[1189]),
      .f(~input_layer[1530]),
      .y(Y[557]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron558_1
  function_37 neuron558_1 (
      .a(input_layer[828]),
      .b(input_layer[1003]),
      .c(~input_layer[1205]),
      .d(input_layer[1259]),
      .e(input_layer[1234]),
      .f(input_layer[1287]),
      .y(Y[558]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron559_1
  function_3 neuron559_1 (
      .a(~input_layer[1429]),
      .b(~input_layer[77]),
      .c(~input_layer[1434]),
      .d(~input_layer[1105]),
      .y(Y[559]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron560_1
  function_42 neuron560_1 (
      .a(input_layer[1219]),
      .b(input_layer[569]),
      .c(input_layer[1280]),
      .d(~input_layer[814]),
      .y(Y[560]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron561_1
  function_27 neuron561_1 (
      .a(~input_layer[967]),
      .b(~input_layer[962]),
      .c(input_layer[1035]),
      .y(Y[561]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron562_1
  function_47 neuron562_1 (
      .a(input_layer[940]),
      .b(input_layer[463]),
      .c(input_layer[190]),
      .d(input_layer[750]),
      .e(input_layer[1312]),
      .y(Y[562]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_209 for neuron563_1
  function_209 neuron563_1 (
      .a(~input_layer[384]),
      .b(input_layer[1539]),
      .c(input_layer[244]),
      .d(input_layer[1359]),
      .e(input_layer[948]),
      .f(input_layer[395]),
      .y(Y[563]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron564_1
  function_35 neuron564_1 (
      .a(~input_layer[1133]),
      .b(~input_layer[756]),
      .c(~input_layer[363]),
      .d(input_layer[927]),
      .e(~input_layer[1395]),
      .y(Y[564]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron565_1
  function_172 neuron565_1 (
      .a(~input_layer[548]),
      .b(~input_layer[1081]),
      .c(~input_layer[919]),
      .d(~input_layer[452]),
      .e(input_layer[1035]),
      .f(~input_layer[667]),
      .y(Y[565]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron566_1
  function_48 neuron566_1 (
      .a(input_layer[680]),
      .b(input_layer[1186]),
      .c(input_layer[1245]),
      .d(~input_layer[270]),
      .e(input_layer[892]),
      .y(Y[566]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron567_1
  function_210 neuron567_1 (
      .a(input_layer[554]),
      .b(~input_layer[143]),
      .c(~input_layer[1125]),
      .d(~input_layer[1468]),
      .e(~input_layer[1472]),
      .f(~input_layer[1435]),
      .y(Y[567]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron568_1
  function_35 neuron568_1 (
      .a(~input_layer[253]),
      .b(input_layer[690]),
      .c(~input_layer[306]),
      .d(~input_layer[1075]),
      .e(~input_layer[130]),
      .y(Y[568]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron569_1
  function_42 neuron569_1 (
      .a(input_layer[460]),
      .b(input_layer[1438]),
      .c(~input_layer[592]),
      .d(input_layer[333]),
      .y(Y[569]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron570_1
  function_24 neuron570_1 (
      .a(~input_layer[1035]),
      .b(~input_layer[322]),
      .c(input_layer[1294]),
      .y(Y[570]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_211 for neuron571_1
  function_211 neuron571_1 (
      .a(~input_layer[387]),
      .b(~input_layer[1022]),
      .c(input_layer[1486]),
      .d(~input_layer[414]),
      .e(input_layer[676]),
      .f(input_layer[673]),
      .y(Y[571]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron572_1
  function_93 neuron572_1 (
      .a(~input_layer[591]),
      .b(input_layer[154]),
      .c(input_layer[864]),
      .d(~input_layer[484]),
      .e(~input_layer[341]),
      .y(Y[572]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron573_1
  function_146 neuron573_1 (
      .a(input_layer[488]),
      .b(input_layer[706]),
      .c(input_layer[149]),
      .d(~input_layer[758]),
      .e(input_layer[1434]),
      .f(~input_layer[286]),
      .y(Y[573]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron574_1
  function_90 neuron574_1 (
      .a(~input_layer[429]),
      .b(input_layer[1091]),
      .c(~input_layer[289]),
      .d(~input_layer[470]),
      .e(input_layer[96]),
      .y(Y[574]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_212 for neuron575_1
  function_212 neuron575_1 (
      .a(input_layer[629]),
      .b(input_layer[795]),
      .c(~input_layer[1334]),
      .d(~input_layer[850]),
      .e(input_layer[670]),
      .y(Y[575]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_213 for neuron576_1
  function_213 neuron576_1 (
      .a(input_layer[1494]),
      .b(input_layer[930]),
      .c(~input_layer[1115]),
      .d(~input_layer[1151]),
      .e(~input_layer[1055]),
      .f(input_layer[1094]),
      .y(Y[576]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron577_1
  function_126 neuron577_1 (
      .a(~input_layer[1296]),
      .b(~input_layer[1077]),
      .c(input_layer[879]),
      .d(~input_layer[550]),
      .e(~input_layer[1471]),
      .y(Y[577]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron578_1
  function_214 neuron578_1 (
      .a(input_layer[1549]),
      .b(input_layer[91]),
      .c(~input_layer[1130]),
      .d(input_layer[96]),
      .e(input_layer[1418]),
      .f(~input_layer[519]),
      .y(Y[578]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_215 for neuron579_1
  function_215 neuron579_1 (
      .a(input_layer[1370]),
      .b(~input_layer[1044]),
      .c(~input_layer[1338]),
      .d(~input_layer[351]),
      .e(~input_layer[123]),
      .f(~input_layer[843]),
      .y(Y[579]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_204 for neuron580_1
  function_204 neuron580_1 (
      .a(~input_layer[1156]),
      .b(input_layer[452]),
      .c(~input_layer[1029]),
      .d(~input_layer[693]),
      .e(input_layer[92]),
      .f(~input_layer[839]),
      .y(Y[580]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron581_1
  function_8 neuron581_1 (
      .a(input_layer[1370]),
      .b(input_layer[1183]),
      .c(input_layer[419]),
      .d(~input_layer[576]),
      .y(Y[581]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron582_1
  function_29 neuron582_1 (
      .a(~input_layer[522]),
      .b(~input_layer[509]),
      .y(Y[582]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron583_1
  function_107 neuron583_1 (
      .a(~input_layer[1017]),
      .b(~input_layer[360]),
      .c(input_layer[126]),
      .d(~input_layer[536]),
      .e(input_layer[507]),
      .y(Y[583]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron584_1
  function_93 neuron584_1 (
      .a(input_layer[189]),
      .b(~input_layer[535]),
      .c(input_layer[195]),
      .d(input_layer[197]),
      .e(~input_layer[589]),
      .y(Y[584]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron585_1
  function_120 neuron585_1 (
      .a(input_layer[715]),
      .b(~input_layer[552]),
      .c(input_layer[596]),
      .d(~input_layer[319]),
      .e(input_layer[779]),
      .y(Y[585]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron586_1
  function_119 neuron586_1 (
      .a(~input_layer[924]),
      .b(~input_layer[1335]),
      .c(~input_layer[782]),
      .d(~input_layer[339]),
      .e(input_layer[1517]),
      .y(Y[586]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron587_1
  function_39 neuron587_1 (
      .a(input_layer[190]),
      .b(input_layer[258]),
      .c(~input_layer[1374]),
      .y(Y[587]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_216 for neuron588_1
  function_216 neuron588_1 (
      .a(input_layer[656]),
      .b(~input_layer[1015]),
      .c(input_layer[622]),
      .d(input_layer[451]),
      .e(~input_layer[1332]),
      .f(input_layer[577]),
      .y(Y[588]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron589_1
  function_31 neuron589_1 (
      .a(~input_layer[1321]),
      .b(input_layer[183]),
      .c(input_layer[766]),
      .d(input_layer[356]),
      .y(Y[589]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron590_1
  function_42 neuron590_1 (
      .a(input_layer[1490]),
      .b(input_layer[1224]),
      .c(input_layer[830]),
      .d(input_layer[1276]),
      .y(Y[590]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_217 for neuron591_1
  function_217 neuron591_1 (
      .a(input_layer[866]),
      .b(~input_layer[424]),
      .c(input_layer[1359]),
      .d(~input_layer[1131]),
      .e(input_layer[1515]),
      .f(input_layer[28]),
      .y(Y[591]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_218 for neuron592_1
  function_218 neuron592_1 (
      .a(input_layer[631]),
      .b(~input_layer[367]),
      .c(input_layer[520]),
      .d(input_layer[1432]),
      .e(~input_layer[1318]),
      .y(Y[592]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_219 for neuron593_1
  function_219 neuron593_1 (
      .a(~input_layer[1190]),
      .b(~input_layer[752]),
      .c(input_layer[651]),
      .d(input_layer[676]),
      .e(input_layer[797]),
      .f(~input_layer[1004]),
      .y(Y[593]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[594] = 1'b0;

  // instantiate function_177 for neuron595_1
  function_177 neuron595_1 (
      .a(~input_layer[1363]),
      .b(~input_layer[1307]),
      .c(input_layer[507]),
      .d(input_layer[430]),
      .e(input_layer[197]),
      .y(Y[595]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_220 for neuron596_1
  function_220 neuron596_1 (
      .a(input_layer[1182]),
      .b(~input_layer[376]),
      .c(~input_layer[434]),
      .d(input_layer[1366]),
      .e(~input_layer[1009]),
      .f(input_layer[26]),
      .y(Y[596]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron597_1
  function_27 neuron597_1 (
      .a(~input_layer[374]),
      .b(~input_layer[1261]),
      .c(~input_layer[1486]),
      .y(Y[597]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron598_1
  function_60 neuron598_1 (
      .a(input_layer[1434]),
      .b(input_layer[1129]),
      .c(~input_layer[420]),
      .d(input_layer[752]),
      .e(~input_layer[942]),
      .y(Y[598]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron599_1
  function_221 neuron599_1 (
      .a(input_layer[1169]),
      .b(~input_layer[1369]),
      .c(input_layer[1152]),
      .d(input_layer[179]),
      .e(input_layer[1154]),
      .f(~input_layer[1513]),
      .y(Y[599]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron600_1
  function_55 neuron600_1 (
      .a(~input_layer[198]),
      .b(~input_layer[1108]),
      .c(input_layer[327]),
      .d(~input_layer[662]),
      .e(~input_layer[276]),
      .y(Y[600]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron601_1
  function_26 neuron601_1 (
      .a(input_layer[1310]),
      .y(Y[601]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron602_1
  function_67 neuron602_1 (
      .a(~input_layer[142]),
      .b(~input_layer[612]),
      .c(~input_layer[565]),
      .d(~input_layer[97]),
      .e(~input_layer[391]),
      .y(Y[602]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron603_1
  function_12 neuron603_1 (
      .a(input_layer[1333]),
      .b(~input_layer[365]),
      .c(input_layer[919]),
      .y(Y[603]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron604_1
  function_97 neuron604_1 (
      .a(~input_layer[764]),
      .b(~input_layer[1385]),
      .c(~input_layer[1384]),
      .d(~input_layer[1391]),
      .e(~input_layer[1043]),
      .y(Y[604]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron605_1
  function_42 neuron605_1 (
      .a(input_layer[1192]),
      .b(input_layer[442]),
      .c(input_layer[703]),
      .d(input_layer[871]),
      .y(Y[605]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron606_1
  function_55 neuron606_1 (
      .a(~input_layer[1138]),
      .b(~input_layer[193]),
      .c(~input_layer[609]),
      .d(input_layer[966]),
      .e(input_layer[1318]),
      .y(Y[606]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_143 for neuron607_1
  function_143 neuron607_1 (
      .a(input_layer[206]),
      .b(input_layer[1494]),
      .c(input_layer[157]),
      .d(~input_layer[552]),
      .e(input_layer[951]),
      .f(input_layer[684]),
      .y(Y[607]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron608_1
  function_17 neuron608_1 (
      .a(input_layer[1053]),
      .b(input_layer[912]),
      .c(~input_layer[645]),
      .y(Y[608]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron609_1
  function_42 neuron609_1 (
      .a(input_layer[1171]),
      .b(input_layer[1546]),
      .c(input_layer[1199]),
      .d(input_layer[1429]),
      .y(Y[609]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron610_1
  function_37 neuron610_1 (
      .a(input_layer[1014]),
      .b(~input_layer[549]),
      .c(input_layer[863]),
      .d(input_layer[233]),
      .e(input_layer[1006]),
      .f(input_layer[1565]),
      .y(Y[610]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_222 for neuron611_1
  function_222 neuron611_1 (
      .a(input_layer[1275]),
      .b(~input_layer[1471]),
      .c(~input_layer[648]),
      .d(input_layer[891]),
      .e(input_layer[1042]),
      .f(input_layer[119]),
      .y(Y[611]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_223 for neuron612_1
  function_223 neuron612_1 (
      .a(input_layer[1426]),
      .b(input_layer[1368]),
      .c(~input_layer[131]),
      .d(input_layer[1302]),
      .e(~input_layer[1223]),
      .f(input_layer[422]),
      .y(Y[612]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_224 for neuron613_1
  function_224 neuron613_1 (
      .a(~input_layer[855]),
      .b(input_layer[463]),
      .c(input_layer[294]),
      .d(~input_layer[131]),
      .e(input_layer[1038]),
      .f(~input_layer[712]),
      .y(Y[613]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_225 for neuron614_1
  function_225 neuron614_1 (
      .a(input_layer[1545]),
      .b(~input_layer[272]),
      .c(input_layer[514]),
      .d(input_layer[654]),
      .e(input_layer[475]),
      .f(input_layer[505]),
      .y(Y[614]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron615_1
  function_181 neuron615_1 (
      .a(~input_layer[1225]),
      .b(input_layer[1540]),
      .c(input_layer[1533]),
      .d(input_layer[674]),
      .e(input_layer[1233]),
      .y(Y[615]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_190 for neuron616_1
  function_190 neuron616_1 (
      .a(~input_layer[1273]),
      .b(input_layer[1540]),
      .c(input_layer[1126]),
      .d(~input_layer[365]),
      .e(~input_layer[1329]),
      .f(input_layer[1061]),
      .y(Y[616]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron617_1
  function_146 neuron617_1 (
      .a(input_layer[441]),
      .b(input_layer[942]),
      .c(input_layer[239]),
      .d(input_layer[946]),
      .e(~input_layer[873]),
      .f(~input_layer[863]),
      .y(Y[617]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron618_1
  function_149 neuron618_1 (
      .a(~input_layer[1369]),
      .b(input_layer[1072]),
      .c(input_layer[1139]),
      .d(~input_layer[1444]),
      .y(Y[618]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron619_1
  function_12 neuron619_1 (
      .a(input_layer[983]),
      .b(~input_layer[1050]),
      .c(input_layer[1165]),
      .y(Y[619]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_226 for neuron620_1
  function_226 neuron620_1 (
      .a(input_layer[931]),
      .b(~input_layer[89]),
      .c(~input_layer[1180]),
      .d(~input_layer[663]),
      .e(~input_layer[662]),
      .f(input_layer[691]),
      .y(Y[620]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_227 for neuron621_1
  function_227 neuron621_1 (
      .a(input_layer[490]),
      .b(~input_layer[244]),
      .c(~input_layer[1348]),
      .d(~input_layer[214]),
      .e(~input_layer[1112]),
      .f(~input_layer[1406]),
      .y(Y[621]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron622_1
  function_12 neuron622_1 (
      .a(input_layer[261]),
      .b(~input_layer[1485]),
      .c(~input_layer[1467]),
      .y(Y[622]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_228 for neuron623_1
  function_228 neuron623_1 (
      .a(input_layer[1202]),
      .b(input_layer[829]),
      .c(~input_layer[329]),
      .d(input_layer[262]),
      .e(input_layer[642]),
      .f(input_layer[664]),
      .y(Y[623]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_229 for neuron624_1
  function_229 neuron624_1 (
      .a(~input_layer[753]),
      .b(~input_layer[661]),
      .c(input_layer[1017]),
      .d(~input_layer[143]),
      .e(~input_layer[666]),
      .f(input_layer[904]),
      .y(Y[624]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron625_1
  function_78 neuron625_1 (
      .a(input_layer[797]),
      .b(~input_layer[890]),
      .c(~input_layer[93]),
      .d(input_layer[1106]),
      .e(~input_layer[842]),
      .f(input_layer[1286]),
      .y(Y[625]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron626_1
  function_157 neuron626_1 (
      .a(input_layer[973]),
      .b(input_layer[372]),
      .c(~input_layer[1407]),
      .d(~input_layer[177]),
      .e(~input_layer[212]),
      .f(input_layer[1453]),
      .y(Y[626]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron627_1
  function_74 neuron627_1 (
      .a(~input_layer[1538]),
      .b(~input_layer[715]),
      .c(~input_layer[1203]),
      .d(~input_layer[1017]),
      .e(input_layer[372]),
      .f(~input_layer[1341]),
      .y(Y[627]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron628_1
  function_27 neuron628_1 (
      .a(~input_layer[1311]),
      .b(~input_layer[1225]),
      .c(input_layer[1142]),
      .y(Y[628]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_230 for neuron629_1
  function_230 neuron629_1 (
      .a(input_layer[500]),
      .b(~input_layer[1482]),
      .c(input_layer[329]),
      .d(input_layer[1318]),
      .e(~input_layer[570]),
      .y(Y[629]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron630_1
  function_29 neuron630_1 (
      .a(~input_layer[807]),
      .b(~input_layer[719]),
      .y(Y[630]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron631_1
  function_39 neuron631_1 (
      .a(input_layer[266]),
      .b(~input_layer[407]),
      .c(~input_layer[1040]),
      .y(Y[631]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron632_1
  function_47 neuron632_1 (
      .a(input_layer[206]),
      .b(input_layer[1168]),
      .c(input_layer[528]),
      .d(input_layer[879]),
      .e(input_layer[947]),
      .y(Y[632]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron633_1
  function_231 neuron633_1 (
      .a(input_layer[837]),
      .b(input_layer[1252]),
      .c(input_layer[1264]),
      .d(input_layer[297]),
      .e(input_layer[390]),
      .f(~input_layer[402]),
      .y(Y[633]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron634_1
  function_26 neuron634_1 (
      .a(input_layer[208]),
      .y(Y[634]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron635_1
  function_232 neuron635_1 (
      .a(~input_layer[983]),
      .b(input_layer[1383]),
      .c(input_layer[1299]),
      .d(~input_layer[237]),
      .e(~input_layer[22]),
      .f(~input_layer[223]),
      .y(Y[635]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron636_1
  function_24 neuron636_1 (
      .a(~input_layer[638]),
      .b(input_layer[1116]),
      .c(input_layer[370]),
      .y(Y[636]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron637_1
  function_67 neuron637_1 (
      .a(~input_layer[1190]),
      .b(~input_layer[1536]),
      .c(~input_layer[945]),
      .d(~input_layer[424]),
      .e(~input_layer[1442]),
      .y(Y[637]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron638_1
  function_29 neuron638_1 (
      .a(~input_layer[377]),
      .b(input_layer[540]),
      .y(Y[638]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron639_1
  function_19 neuron639_1 (
      .a(~input_layer[204]),
      .b(~input_layer[212]),
      .c(~input_layer[129]),
      .d(input_layer[930]),
      .y(Y[639]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron640_1
  function_87 neuron640_1 (
      .a(input_layer[1001]),
      .b(input_layer[1196]),
      .c(~input_layer[1444]),
      .d(input_layer[772]),
      .e(~input_layer[853]),
      .y(Y[640]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron641_1
  function_18 neuron641_1 (
      .a(~input_layer[367]),
      .b(input_layer[1426]),
      .c(~input_layer[1079]),
      .d(~input_layer[777]),
      .e(input_layer[600]),
      .y(Y[641]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron642_1
  function_3 neuron642_1 (
      .a(~input_layer[142]),
      .b(~input_layer[1248]),
      .c(~input_layer[1302]),
      .d(~input_layer[1547]),
      .y(Y[642]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron643_1
  function_30 neuron643_1 (
      .a(input_layer[1079]),
      .b(input_layer[974]),
      .c(~input_layer[1411]),
      .d(input_layer[84]),
      .y(Y[643]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron644_1
  function_167 neuron644_1 (
      .a(input_layer[309]),
      .b(input_layer[389]),
      .c(input_layer[902]),
      .d(~input_layer[766]),
      .e(~input_layer[1374]),
      .y(Y[644]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_233 for neuron645_1
  function_233 neuron645_1 (
      .a(~input_layer[537]),
      .b(input_layer[358]),
      .c(~input_layer[299]),
      .d(~input_layer[781]),
      .e(input_layer[252]),
      .f(~input_layer[61]),
      .y(Y[645]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron646_1
  function_126 neuron646_1 (
      .a(~input_layer[655]),
      .b(~input_layer[1112]),
      .c(input_layer[399]),
      .d(~input_layer[1547]),
      .e(~input_layer[792]),
      .y(Y[646]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron647_1
  function_26 neuron647_1 (
      .a(input_layer[1034]),
      .y(Y[647]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron648_1
  function_67 neuron648_1 (
      .a(~input_layer[290]),
      .b(~input_layer[1092]),
      .c(~input_layer[453]),
      .d(~input_layer[462]),
      .e(~input_layer[781]),
      .y(Y[648]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron649_1
  function_234 neuron649_1 (
      .a(~input_layer[499]),
      .b(~input_layer[383]),
      .c(input_layer[705]),
      .d(~input_layer[213]),
      .e(~input_layer[1557]),
      .f(input_layer[1413]),
      .y(Y[649]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron650_1
  function_25 neuron650_1 (
      .a(~input_layer[476]),
      .b(input_layer[1294]),
      .c(input_layer[1253]),
      .d(input_layer[959]),
      .e(input_layer[974]),
      .y(Y[650]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron651_1
  function_99 neuron651_1 (
      .a(input_layer[1411]),
      .b(input_layer[705]),
      .c(input_layer[959]),
      .d(~input_layer[800]),
      .e(input_layer[1050]),
      .y(Y[651]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron652_1
  function_12 neuron652_1 (
      .a(input_layer[1431]),
      .b(~input_layer[82]),
      .c(input_layer[438]),
      .y(Y[652]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron653_1
  function_48 neuron653_1 (
      .a(input_layer[621]),
      .b(~input_layer[934]),
      .c(input_layer[669]),
      .d(input_layer[387]),
      .e(input_layer[344]),
      .y(Y[653]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_235 for neuron654_1
  function_235 neuron654_1 (
      .a(~input_layer[1429]),
      .b(~input_layer[772]),
      .c(input_layer[1227]),
      .d(~input_layer[383]),
      .e(input_layer[971]),
      .y(Y[654]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_236 for neuron655_1
  function_236 neuron655_1 (
      .a(input_layer[258]),
      .b(~input_layer[874]),
      .c(input_layer[536]),
      .d(input_layer[510]),
      .e(input_layer[605]),
      .f(input_layer[526]),
      .y(Y[655]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_237 for neuron656_1
  function_237 neuron656_1 (
      .a(input_layer[1186]),
      .b(input_layer[454]),
      .c(~input_layer[1117]),
      .d(~input_layer[1548]),
      .e(~input_layer[1382]),
      .y(Y[656]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron657_1
  function_1 neuron657_1 (
      .a(~input_layer[478]),
      .b(~input_layer[454]),
      .c(~input_layer[1536]),
      .d(input_layer[490]),
      .y(Y[657]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron658_1
  function_8 neuron658_1 (
      .a(input_layer[922]),
      .b(input_layer[647]),
      .c(input_layer[333]),
      .d(~input_layer[830]),
      .y(Y[658]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron659_1
  function_55 neuron659_1 (
      .a(~input_layer[936]),
      .b(~input_layer[1280]),
      .c(~input_layer[1467]),
      .d(input_layer[719]),
      .e(~input_layer[391]),
      .y(Y[659]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_238 for neuron660_1
  function_238 neuron660_1 (
      .a(input_layer[329]),
      .b(~input_layer[1189]),
      .c(input_layer[522]),
      .d(~input_layer[566]),
      .e(input_layer[391]),
      .y(Y[660]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_239 for neuron661_1
  function_239 neuron661_1 (
      .a(input_layer[311]),
      .b(~input_layer[819]),
      .c(input_layer[518]),
      .d(input_layer[94]),
      .e(input_layer[1271]),
      .f(input_layer[1292]),
      .y(Y[661]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron662_1
  function_3 neuron662_1 (
      .a(~input_layer[1471]),
      .b(~input_layer[290]),
      .c(~input_layer[1228]),
      .d(~input_layer[819]),
      .y(Y[662]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron663_1
  function_67 neuron663_1 (
      .a(~input_layer[145]),
      .b(~input_layer[721]),
      .c(~input_layer[1542]),
      .d(~input_layer[158]),
      .e(~input_layer[733]),
      .y(Y[663]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron664_1
  function_123 neuron664_1 (
      .a(input_layer[809]),
      .b(~input_layer[1186]),
      .c(~input_layer[1211]),
      .d(input_layer[267]),
      .y(Y[664]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron665_1
  function_7 neuron665_1 (
      .a(input_layer[297]),
      .b(input_layer[548]),
      .c(~input_layer[913]),
      .d(~input_layer[917]),
      .y(Y[665]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron666_1
  function_17 neuron666_1 (
      .a(input_layer[385]),
      .b(input_layer[471]),
      .c(input_layer[82]),
      .y(Y[666]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_240 for neuron667_1
  function_240 neuron667_1 (
      .a(~input_layer[1318]),
      .b(input_layer[978]),
      .c(input_layer[1443]),
      .d(input_layer[1146]),
      .e(~input_layer[598]),
      .f(input_layer[771]),
      .y(Y[667]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron668_1
  function_3 neuron668_1 (
      .a(~input_layer[1486]),
      .b(~input_layer[1169]),
      .c(input_layer[1258]),
      .d(~input_layer[1273]),
      .y(Y[668]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron669_1
  function_241 neuron669_1 (
      .a(input_layer[909]),
      .b(input_layer[1538]),
      .c(input_layer[833]),
      .d(input_layer[1358]),
      .e(input_layer[1431]),
      .f(~input_layer[1387]),
      .y(Y[669]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron670_1
  function_48 neuron670_1 (
      .a(input_layer[1539]),
      .b(input_layer[243]),
      .c(input_layer[159]),
      .d(~input_layer[319]),
      .e(input_layer[216]),
      .y(Y[670]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron671_1
  function_242 neuron671_1 (
      .a(~input_layer[661]),
      .b(input_layer[1181]),
      .c(input_layer[96]),
      .d(~input_layer[833]),
      .e(input_layer[559]),
      .f(~input_layer[590]),
      .y(Y[671]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron672_1
  function_3 neuron672_1 (
      .a(~input_layer[769]),
      .b(~input_layer[1469]),
      .c(~input_layer[261]),
      .d(input_layer[1133]),
      .y(Y[672]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron673_1
  function_27 neuron673_1 (
      .a(~input_layer[750]),
      .b(~input_layer[1044]),
      .c(~input_layer[1076]),
      .y(Y[673]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron674_1
  function_3 neuron674_1 (
      .a(~input_layer[1115]),
      .b(~input_layer[987]),
      .c(~input_layer[957]),
      .d(input_layer[1550]),
      .y(Y[674]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_243 for neuron675_1
  function_243 neuron675_1 (
      .a(~input_layer[741]),
      .b(input_layer[403]),
      .c(input_layer[775]),
      .d(input_layer[675]),
      .e(~input_layer[985]),
      .f(~input_layer[632]),
      .y(Y[675]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron676_1
  function_67 neuron676_1 (
      .a(~input_layer[1014]),
      .b(~input_layer[1478]),
      .c(~input_layer[1005]),
      .d(~input_layer[1069]),
      .e(~input_layer[740]),
      .y(Y[676]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_244 for neuron677_1
  function_244 neuron677_1 (
      .a(~input_layer[1353]),
      .b(input_layer[917]),
      .c(input_layer[1493]),
      .d(~input_layer[288]),
      .e(input_layer[617]),
      .f(input_layer[505]),
      .y(Y[677]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_245 for neuron678_1
  function_245 neuron678_1 (
      .a(input_layer[625]),
      .b(~input_layer[263]),
      .c(~input_layer[1144]),
      .d(~input_layer[684]),
      .e(input_layer[1063]),
      .f(~input_layer[1515]),
      .y(Y[678]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron679_1
  function_202 neuron679_1 (
      .a(~input_layer[1126]),
      .b(~input_layer[1298]),
      .c(~input_layer[1353]),
      .d(input_layer[668]),
      .e(input_layer[871]),
      .f(~input_layer[1272]),
      .y(Y[679]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron680_1
  function_35 neuron680_1 (
      .a(~input_layer[1050]),
      .b(~input_layer[1303]),
      .c(input_layer[810]),
      .d(input_layer[761]),
      .e(~input_layer[1319]),
      .y(Y[680]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron681_1
  function_7 neuron681_1 (
      .a(input_layer[1158]),
      .b(input_layer[1255]),
      .c(~input_layer[143]),
      .d(input_layer[131]),
      .y(Y[681]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron682_1
  function_214 neuron682_1 (
      .a(input_layer[767]),
      .b(input_layer[126]),
      .c(~input_layer[267]),
      .d(~input_layer[926]),
      .e(input_layer[1452]),
      .f(input_layer[70]),
      .y(Y[682]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron683_1
  function_214 neuron683_1 (
      .a(input_layer[766]),
      .b(input_layer[400]),
      .c(input_layer[1182]),
      .d(~input_layer[863]),
      .e(input_layer[1381]),
      .f(~input_layer[1418]),
      .y(Y[683]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron684_1
  function_92 neuron684_1 (
      .a(input_layer[199]),
      .b(input_layer[203]),
      .c(input_layer[1161]),
      .d(input_layer[1115]),
      .e(input_layer[1086]),
      .f(~input_layer[407]),
      .y(Y[684]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_166 for neuron685_1
  function_166 neuron685_1 (
      .a(~input_layer[692]),
      .b(input_layer[644]),
      .c(input_layer[1214]),
      .d(input_layer[1320]),
      .e(input_layer[176]),
      .f(input_layer[119]),
      .y(Y[685]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron686_1
  function_123 neuron686_1 (
      .a(input_layer[1022]),
      .b(~input_layer[453]),
      .c(input_layer[1253]),
      .d(~input_layer[489]),
      .y(Y[686]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_246 for neuron687_1
  function_246 neuron687_1 (
      .a(~input_layer[1242]),
      .b(input_layer[1004]),
      .c(~input_layer[458]),
      .d(input_layer[1440]),
      .e(~input_layer[1192]),
      .f(input_layer[375]),
      .y(Y[687]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_247 for neuron688_1
  function_247 neuron688_1 (
      .a(input_layer[1109]),
      .b(input_layer[859]),
      .c(input_layer[201]),
      .d(~input_layer[1080]),
      .e(input_layer[834]),
      .f(~input_layer[489]),
      .y(Y[688]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron689_1
  function_155 neuron689_1 (
      .a(~input_layer[147]),
      .b(~input_layer[1410]),
      .c(input_layer[1251]),
      .d(input_layer[1134]),
      .e(~input_layer[1145]),
      .f(~input_layer[1406]),
      .y(Y[689]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron690_1
  function_35 neuron690_1 (
      .a(~input_layer[1494]),
      .b(input_layer[870]),
      .c(input_layer[868]),
      .d(~input_layer[1060]),
      .e(input_layer[749]),
      .y(Y[690]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron691_1
  function_42 neuron691_1 (
      .a(input_layer[709]),
      .b(input_layer[1383]),
      .c(input_layer[158]),
      .d(input_layer[610]),
      .y(Y[691]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron692_1
  function_67 neuron692_1 (
      .a(~input_layer[1477]),
      .b(~input_layer[1368]),
      .c(~input_layer[1205]),
      .d(~input_layer[703]),
      .e(~input_layer[834]),
      .y(Y[692]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron693_1
  function_27 neuron693_1 (
      .a(~input_layer[935]),
      .b(~input_layer[1418]),
      .c(~input_layer[1219]),
      .y(Y[693]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron694_1
  function_7 neuron694_1 (
      .a(~input_layer[254]),
      .b(input_layer[667]),
      .c(~input_layer[661]),
      .d(~input_layer[1249]),
      .y(Y[694]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron695_1
  function_120 neuron695_1 (
      .a(input_layer[741]),
      .b(input_layer[745]),
      .c(~input_layer[76]),
      .d(~input_layer[108]),
      .e(~input_layer[839]),
      .y(Y[695]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron696_1
  function_75 neuron696_1 (
      .a(input_layer[1497]),
      .b(~input_layer[907]),
      .c(~input_layer[331]),
      .d(input_layer[237]),
      .e(input_layer[1551]),
      .y(Y[696]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron697_1
  function_248 neuron697_1 (
      .a(~input_layer[701]),
      .b(~input_layer[388]),
      .c(input_layer[659]),
      .d(input_layer[536]),
      .e(input_layer[933]),
      .f(input_layer[1387]),
      .y(Y[697]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron698_1
  function_0 neuron698_1 (
      .a(~input_layer[317]),
      .b(~input_layer[611]),
      .c(~input_layer[607]),
      .d(~input_layer[430]),
      .e(input_layer[819]),
      .y(Y[698]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron699_1
  function_8 neuron699_1 (
      .a(input_layer[1071]),
      .b(input_layer[513]),
      .c(~input_layer[777]),
      .d(~input_layer[1134]),
      .y(Y[699]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron700_1
  function_27 neuron700_1 (
      .a(~input_layer[1484]),
      .b(~input_layer[1478]),
      .c(~input_layer[1422]),
      .y(Y[700]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_237 for neuron701_1
  function_237 neuron701_1 (
      .a(input_layer[382]),
      .b(input_layer[520]),
      .c(~input_layer[77]),
      .d(~input_layer[1045]),
      .e(~input_layer[1348]),
      .y(Y[701]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron702_1
  function_27 neuron702_1 (
      .a(input_layer[1090]),
      .b(~input_layer[130]),
      .c(~input_layer[1199]),
      .y(Y[702]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_249 for neuron703_1
  function_249 neuron703_1 (
      .a(~input_layer[750]),
      .b(~input_layer[245]),
      .c(~input_layer[855]),
      .d(input_layer[1538]),
      .e(input_layer[397]),
      .y(Y[703]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron704_1
  function_148 neuron704_1 (
      .a(input_layer[777]),
      .b(input_layer[1283]),
      .c(input_layer[1151]),
      .d(~input_layer[192]),
      .e(input_layer[783]),
      .f(~input_layer[952]),
      .y(Y[704]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_250 for neuron705_1
  function_250 neuron705_1 (
      .a(~input_layer[1217]),
      .b(input_layer[1447]),
      .c(~input_layer[412]),
      .d(~input_layer[1303]),
      .e(input_layer[1232]),
      .f(input_layer[1505]),
      .y(Y[705]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron706_1
  function_123 neuron706_1 (
      .a(input_layer[1492]),
      .b(~input_layer[704]),
      .c(~input_layer[353]),
      .d(~input_layer[734]),
      .y(Y[706]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron707_1
  function_242 neuron707_1 (
      .a(input_layer[1438]),
      .b(input_layer[1470]),
      .c(~input_layer[940]),
      .d(input_layer[712]),
      .e(~input_layer[1038]),
      .f(input_layer[390]),
      .y(Y[707]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron708_1
  function_1 neuron708_1 (
      .a(~input_layer[500]),
      .b(input_layer[1206]),
      .c(~input_layer[197]),
      .d(~input_layer[709]),
      .y(Y[708]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron709_1
  function_26 neuron709_1 (
      .a(~input_layer[855]),
      .y(Y[709]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron710_1
  function_29 neuron710_1 (
      .a(~input_layer[1138]),
      .b(~input_layer[1057]),
      .y(Y[710]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron711_1
  function_12 neuron711_1 (
      .a(~input_layer[550]),
      .b(input_layer[1071]),
      .c(input_layer[966]),
      .y(Y[711]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron712_1
  function_42 neuron712_1 (
      .a(input_layer[202]),
      .b(input_layer[781]),
      .c(input_layer[89]),
      .d(~input_layer[1205]),
      .y(Y[712]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron713_1
  function_99 neuron713_1 (
      .a(input_layer[891]),
      .b(input_layer[1087]),
      .c(~input_layer[609]),
      .d(input_layer[1015]),
      .e(input_layer[1529]),
      .y(Y[713]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron714_1
  function_12 neuron714_1 (
      .a(input_layer[922]),
      .b(~input_layer[969]),
      .c(input_layer[1357]),
      .y(Y[714]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_251 for neuron715_1
  function_251 neuron715_1 (
      .a(input_layer[1136]),
      .b(input_layer[1245]),
      .c(~input_layer[1432]),
      .d(~input_layer[741]),
      .e(input_layer[855]),
      .f(~input_layer[671]),
      .y(Y[715]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_252 for neuron716_1
  function_252 neuron716_1 (
      .a(~input_layer[492]),
      .b(input_layer[142]),
      .c(~input_layer[1258]),
      .d(~input_layer[1249]),
      .e(~input_layer[855]),
      .f(input_layer[1556]),
      .y(Y[716]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron717_1
  function_29 neuron717_1 (
      .a(~input_layer[314]),
      .b(~input_layer[411]),
      .y(Y[717]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron718_1
  function_36 neuron718_1 (
      .a(input_layer[242]),
      .b(input_layer[1124]),
      .c(input_layer[90]),
      .d(~input_layer[467]),
      .e(input_layer[1382]),
      .f(~input_layer[1409]),
      .y(Y[718]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron719_1
  function_12 neuron719_1 (
      .a(input_layer[437]),
      .b(input_layer[208]),
      .c(~input_layer[1490]),
      .y(Y[719]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron720_1
  function_4 neuron720_1 (
      .a(~input_layer[972]),
      .b(~input_layer[974]),
      .c(~input_layer[620]),
      .d(input_layer[1134]),
      .e(~input_layer[269]),
      .y(Y[720]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron721_1
  function_27 neuron721_1 (
      .a(input_layer[1136]),
      .b(~input_layer[1436]),
      .c(~input_layer[1496]),
      .y(Y[721]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron722_1
  function_155 neuron722_1 (
      .a(~input_layer[202]),
      .b(~input_layer[883]),
      .c(~input_layer[1171]),
      .d(~input_layer[1539]),
      .e(~input_layer[602]),
      .f(input_layer[529]),
      .y(Y[722]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron723_1
  function_29 neuron723_1 (
      .a(~input_layer[1071]),
      .b(input_layer[1137]),
      .y(Y[723]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron724_1
  function_11 neuron724_1 (
      .a(~input_layer[983]),
      .b(input_layer[472]),
      .c(~input_layer[1128]),
      .d(input_layer[996]),
      .y(Y[724]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron725_1
  function_186 neuron725_1 (
      .a(input_layer[1274]),
      .b(input_layer[1435]),
      .c(~input_layer[943]),
      .d(~input_layer[91]),
      .y(Y[725]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron726_1
  function_253 neuron726_1 (
      .a(input_layer[979]),
      .b(input_layer[498]),
      .c(input_layer[1303]),
      .d(input_layer[1198]),
      .e(~input_layer[1548]),
      .f(input_layer[295]),
      .y(Y[726]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_254 for neuron727_1
  function_254 neuron727_1 (
      .a(~input_layer[388]),
      .b(~input_layer[323]),
      .c(~input_layer[308]),
      .d(input_layer[521]),
      .e(input_layer[607]),
      .f(input_layer[1381]),
      .y(Y[727]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron728_1
  function_30 neuron728_1 (
      .a(input_layer[1326]),
      .b(input_layer[1248]),
      .c(input_layer[620]),
      .d(~input_layer[856]),
      .y(Y[728]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron729_1
  function_42 neuron729_1 (
      .a(input_layer[142]),
      .b(input_layer[644]),
      .c(input_layer[514]),
      .d(input_layer[343]),
      .y(Y[729]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron730_1
  function_74 neuron730_1 (
      .a(input_layer[716]),
      .b(~input_layer[1181]),
      .c(~input_layer[724]),
      .d(~input_layer[1041]),
      .e(~input_layer[162]),
      .f(~input_layer[822]),
      .y(Y[730]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron731_1
  function_5 neuron731_1 (
      .a(~input_layer[991]),
      .b(~input_layer[1296]),
      .c(~input_layer[288]),
      .d(~input_layer[1553]),
      .e(input_layer[269]),
      .f(input_layer[436]),
      .y(Y[731]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron732_1
  function_42 neuron732_1 (
      .a(input_layer[1020]),
      .b(input_layer[1048]),
      .c(input_layer[1154]),
      .d(input_layer[999]),
      .y(Y[732]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron733_1
  function_27 neuron733_1 (
      .a(~input_layer[917]),
      .b(~input_layer[1141]),
      .c(~input_layer[1169]),
      .y(Y[733]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron734_1
  function_27 neuron734_1 (
      .a(~input_layer[349]),
      .b(~input_layer[763]),
      .c(input_layer[316]),
      .y(Y[734]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron735_1
  function_97 neuron735_1 (
      .a(~input_layer[540]),
      .b(input_layer[1026]),
      .c(~input_layer[464]),
      .d(~input_layer[1530]),
      .e(~input_layer[1448]),
      .y(Y[735]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron736_1
  function_56 neuron736_1 (
      .a(~input_layer[803]),
      .b(input_layer[1544]),
      .c(input_layer[1091]),
      .d(input_layer[724]),
      .e(~input_layer[1265]),
      .y(Y[736]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron737_1
  function_52 neuron737_1 (
      .a(~input_layer[1112]),
      .b(input_layer[530]),
      .c(input_layer[509]),
      .d(input_layer[248]),
      .e(input_layer[1357]),
      .f(input_layer[27]),
      .y(Y[737]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron738_1
  function_78 neuron738_1 (
      .a(~input_layer[746]),
      .b(~input_layer[794]),
      .c(~input_layer[139]),
      .d(~input_layer[1192]),
      .e(~input_layer[1237]),
      .f(input_layer[58]),
      .y(Y[738]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_255 for neuron739_1
  function_255 neuron739_1 (
      .a(~input_layer[902]),
      .b(input_layer[1031]),
      .c(input_layer[747]),
      .d(~input_layer[926]),
      .e(input_layer[1205]),
      .y(Y[739]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron740_1
  function_26 neuron740_1 (
      .a(input_layer[1018]),
      .y(Y[740]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[741] = 1'b1;

  // instantiate function_107 for neuron742_1
  function_107 neuron742_1 (
      .a(input_layer[753]),
      .b(~input_layer[237]),
      .c(~input_layer[452]),
      .d(~input_layer[618]),
      .e(input_layer[125]),
      .y(Y[742]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron743_1
  function_30 neuron743_1 (
      .a(input_layer[907]),
      .b(input_layer[1335]),
      .c(~input_layer[1499]),
      .d(~input_layer[74]),
      .y(Y[743]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_256 for neuron744_1
  function_256 neuron744_1 (
      .a(input_layer[776]),
      .b(input_layer[639]),
      .c(input_layer[136]),
      .d(~input_layer[239]),
      .e(input_layer[1085]),
      .f(~input_layer[649]),
      .y(Y[744]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_15 for neuron745_1
  function_15 neuron745_1 (
      .a(input_layer[687]),
      .b(input_layer[582]),
      .c(~input_layer[650]),
      .d(input_layer[525]),
      .e(input_layer[883]),
      .f(input_layer[766]),
      .y(Y[745]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_257 for neuron746_1
  function_257 neuron746_1 (
      .a(input_layer[525]),
      .b(input_layer[87]),
      .c(input_layer[710]),
      .d(input_layer[532]),
      .e(~input_layer[968]),
      .f(input_layer[1356]),
      .y(Y[746]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron747_1
  function_24 neuron747_1 (
      .a(~input_layer[911]),
      .b(input_layer[669]),
      .c(~input_layer[485]),
      .y(Y[747]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron748_1
  function_16 neuron748_1 (
      .a(input_layer[660]),
      .b(input_layer[712]),
      .y(Y[748]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron749_1
  function_8 neuron749_1 (
      .a(input_layer[860]),
      .b(input_layer[968]),
      .c(input_layer[131]),
      .d(~input_layer[1472]),
      .y(Y[749]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron750_1
  function_17 neuron750_1 (
      .a(input_layer[827]),
      .b(input_layer[824]),
      .c(input_layer[1072]),
      .y(Y[750]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron751_1
  function_17 neuron751_1 (
      .a(input_layer[346]),
      .b(input_layer[243]),
      .c(input_layer[209]),
      .y(Y[751]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_258 for neuron752_1
  function_258 neuron752_1 (
      .a(~input_layer[237]),
      .b(input_layer[854]),
      .c(input_layer[1494]),
      .d(~input_layer[1083]),
      .e(~input_layer[1028]),
      .f(input_layer[791]),
      .y(Y[752]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_259 for neuron753_1
  function_259 neuron753_1 (
      .a(~input_layer[1440]),
      .b(input_layer[594]),
      .c(input_layer[396]),
      .d(input_layer[516]),
      .e(~input_layer[603]),
      .y(Y[753]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[754] = 1'b1;

  // instantiate function_8 for neuron755_1
  function_8 neuron755_1 (
      .a(input_layer[1280]),
      .b(input_layer[349]),
      .c(~input_layer[807]),
      .d(~input_layer[311]),
      .y(Y[755]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron756_1
  function_26 neuron756_1 (
      .a(~input_layer[750]),
      .y(Y[756]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_260 for neuron757_1
  function_260 neuron757_1 (
      .a(~input_layer[773]),
      .b(~input_layer[1365]),
      .c(input_layer[1297]),
      .d(input_layer[900]),
      .e(~input_layer[1303]),
      .f(input_layer[794]),
      .y(Y[757]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_261 for neuron758_1
  function_261 neuron758_1 (
      .a(input_layer[816]),
      .b(~input_layer[1109]),
      .c(~input_layer[1253]),
      .d(input_layer[557]),
      .e(input_layer[287]),
      .f(~input_layer[1092]),
      .y(Y[758]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[759] = 1'b0;

  // instantiate function_262 for neuron760_1
  function_262 neuron760_1 (
      .a(input_layer[772]),
      .b(input_layer[889]),
      .c(~input_layer[1294]),
      .d(input_layer[1155]),
      .e(~input_layer[437]),
      .f(~input_layer[685]),
      .y(Y[760]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron761_1
  function_7 neuron761_1 (
      .a(input_layer[1241]),
      .b(input_layer[484]),
      .c(~input_layer[721]),
      .d(~input_layer[971]),
      .y(Y[761]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron762_1
  function_0 neuron762_1 (
      .a(~input_layer[499]),
      .b(~input_layer[832]),
      .c(~input_layer[93]),
      .d(~input_layer[614]),
      .e(~input_layer[350]),
      .y(Y[762]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron763_1
  function_39 neuron763_1 (
      .a(input_layer[1278]),
      .b(~input_layer[310]),
      .c(~input_layer[1069]),
      .y(Y[763]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron764_1
  function_106 neuron764_1 (
      .a(~input_layer[1237]),
      .b(input_layer[437]),
      .c(input_layer[1132]),
      .d(input_layer[1079]),
      .y(Y[764]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_263 for neuron765_1
  function_263 neuron765_1 (
      .a(~input_layer[260]),
      .b(~input_layer[865]),
      .c(input_layer[408]),
      .d(input_layer[589]),
      .e(input_layer[397]),
      .f(~input_layer[899]),
      .y(Y[765]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_264 for neuron766_1
  function_264 neuron766_1 (
      .a(~input_layer[908]),
      .b(input_layer[146]),
      .c(input_layer[1017]),
      .d(~input_layer[259]),
      .e(~input_layer[1225]),
      .f(~input_layer[1226]),
      .y(Y[766]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_159 for neuron767_1
  function_159 neuron767_1 (
      .a(~input_layer[920]),
      .b(input_layer[255]),
      .c(~input_layer[1041]),
      .d(input_layer[516]),
      .e(input_layer[901]),
      .f(~input_layer[1275]),
      .y(Y[767]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_265 for neuron768_1
  function_265 neuron768_1 (
      .a(~input_layer[347]),
      .b(input_layer[798]),
      .c(input_layer[968]),
      .d(~input_layer[1362]),
      .e(input_layer[641]),
      .f(input_layer[1406]),
      .y(Y[768]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron769_1
  function_67 neuron769_1 (
      .a(~input_layer[261]),
      .b(~input_layer[889]),
      .c(~input_layer[1547]),
      .d(~input_layer[949]),
      .e(~input_layer[92]),
      .y(Y[769]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_266 for neuron770_1
  function_266 neuron770_1 (
      .a(~input_layer[716]),
      .b(input_layer[442]),
      .c(~input_layer[406]),
      .d(input_layer[323]),
      .e(~input_layer[217]),
      .f(~input_layer[883]),
      .y(Y[770]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron771_1
  function_26 neuron771_1 (
      .a(~input_layer[988]),
      .y(Y[771]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_267 for neuron772_1
  function_267 neuron772_1 (
      .a(~input_layer[314]),
      .b(~input_layer[435]),
      .c(~input_layer[669]),
      .d(input_layer[792]),
      .e(input_layer[1302]),
      .f(input_layer[813]),
      .y(Y[772]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_268 for neuron773_1
  function_268 neuron773_1 (
      .a(input_layer[1377]),
      .b(~input_layer[1549]),
      .c(~input_layer[589]),
      .d(~input_layer[732]),
      .e(~input_layer[541]),
      .f(~input_layer[1063]),
      .y(Y[773]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron774_1
  function_27 neuron774_1 (
      .a(input_layer[968]),
      .b(input_layer[1252]),
      .c(input_layer[803]),
      .y(Y[774]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron775_1
  function_120 neuron775_1 (
      .a(~input_layer[384]),
      .b(input_layer[1001]),
      .c(input_layer[298]),
      .d(input_layer[1066]),
      .e(~input_layer[922]),
      .y(Y[775]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_269 for neuron776_1
  function_269 neuron776_1 (
      .a(input_layer[569]),
      .b(input_layer[790]),
      .c(input_layer[788]),
      .d(input_layer[447]),
      .e(input_layer[70]),
      .f(~input_layer[1320]),
      .y(Y[776]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_270 for neuron777_1
  function_270 neuron777_1 (
      .a(input_layer[137]),
      .b(~input_layer[753]),
      .c(input_layer[1356]),
      .d(~input_layer[1336]),
      .e(~input_layer[1312]),
      .f(~input_layer[1209]),
      .y(Y[777]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron778_1
  function_29 neuron778_1 (
      .a(~input_layer[661]),
      .b(~input_layer[1311]),
      .y(Y[778]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron779_1
  function_16 neuron779_1 (
      .a(input_layer[203]),
      .b(~input_layer[426]),
      .y(Y[779]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron780_1
  function_48 neuron780_1 (
      .a(input_layer[611]),
      .b(~input_layer[1142]),
      .c(input_layer[208]),
      .d(input_layer[1528]),
      .e(input_layer[1294]),
      .y(Y[780]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron781_1
  function_29 neuron781_1 (
      .a(~input_layer[1414]),
      .b(~input_layer[822]),
      .y(Y[781]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron782_1
  function_106 neuron782_1 (
      .a(input_layer[1080]),
      .b(input_layer[1543]),
      .c(~input_layer[799]),
      .d(~input_layer[1384]),
      .y(Y[782]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron783_1
  function_47 neuron783_1 (
      .a(input_layer[977]),
      .b(input_layer[1483]),
      .c(input_layer[595]),
      .d(input_layer[949]),
      .e(input_layer[1060]),
      .y(Y[783]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron784_1
  function_48 neuron784_1 (
      .a(input_layer[135]),
      .b(input_layer[1355]),
      .c(~input_layer[925]),
      .d(input_layer[124]),
      .e(input_layer[1090]),
      .y(Y[784]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron785_1
  function_26 neuron785_1 (
      .a(~input_layer[1086]),
      .y(Y[785]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron786_1
  function_7 neuron786_1 (
      .a(input_layer[755]),
      .b(~input_layer[539]),
      .c(input_layer[862]),
      .d(input_layer[863]),
      .y(Y[786]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron787_1
  function_39 neuron787_1 (
      .a(input_layer[498]),
      .b(~input_layer[941]),
      .c(input_layer[1365]),
      .y(Y[787]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron788_1
  function_46 neuron788_1 (
      .a(input_layer[154]),
      .b(input_layer[1541]),
      .c(input_layer[244]),
      .d(~input_layer[1331]),
      .e(~input_layer[428]),
      .y(Y[788]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron789_1
  function_126 neuron789_1 (
      .a(~input_layer[662]),
      .b(~input_layer[187]),
      .c(~input_layer[722]),
      .d(input_layer[1413]),
      .e(~input_layer[1181]),
      .y(Y[789]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron790_1
  function_26 neuron790_1 (
      .a(input_layer[760]),
      .y(Y[790]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron791_1
  function_27 neuron791_1 (
      .a(~input_layer[323]),
      .b(~input_layer[261]),
      .c(~input_layer[495]),
      .y(Y[791]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron792_1
  function_70 neuron792_1 (
      .a(~input_layer[886]),
      .b(~input_layer[241]),
      .c(~input_layer[903]),
      .d(input_layer[414]),
      .e(input_layer[399]),
      .f(input_layer[52]),
      .y(Y[792]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron793_1
  function_17 neuron793_1 (
      .a(input_layer[1017]),
      .b(input_layer[347]),
      .c(input_layer[861]),
      .y(Y[793]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron794_1
  function_26 neuron794_1 (
      .a(~input_layer[977]),
      .y(Y[794]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron795_1
  function_271 neuron795_1 (
      .a(input_layer[188]),
      .b(input_layer[83]),
      .c(input_layer[1203]),
      .d(~input_layer[836]),
      .e(input_layer[1042]),
      .y(Y[795]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron796_1
  function_35 neuron796_1 (
      .a(~input_layer[301]),
      .b(~input_layer[413]),
      .c(~input_layer[544]),
      .d(input_layer[1446]),
      .e(~input_layer[499]),
      .y(Y[796]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron797_1
  function_39 neuron797_1 (
      .a(input_layer[1497]),
      .b(~input_layer[1263]),
      .c(~input_layer[1309]),
      .y(Y[797]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron798_1
  function_30 neuron798_1 (
      .a(input_layer[1199]),
      .b(input_layer[87]),
      .c(input_layer[1108]),
      .d(~input_layer[738]),
      .y(Y[798]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_272 for neuron799_1
  function_272 neuron799_1 (
      .a(input_layer[792]),
      .b(~input_layer[883]),
      .c(~input_layer[159]),
      .d(~input_layer[1316]),
      .e(input_layer[635]),
      .f(input_layer[921]),
      .y(Y[799]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron800_1
  function_67 neuron800_1 (
      .a(~input_layer[344]),
      .b(input_layer[750]),
      .c(~input_layer[1351]),
      .d(~input_layer[241]),
      .e(~input_layer[1529]),
      .y(Y[800]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron801_1
  function_28 neuron801_1 (
      .a(~input_layer[552]),
      .b(~input_layer[1294]),
      .c(~input_layer[400]),
      .d(~input_layer[523]),
      .e(~input_layer[1532]),
      .f(input_layer[988]),
      .y(Y[801]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_273 for neuron802_1
  function_273 neuron802_1 (
      .a(~input_layer[1417]),
      .b(input_layer[1164]),
      .c(input_layer[1078]),
      .d(~input_layer[401]),
      .e(input_layer[1173]),
      .y(Y[802]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[803] = 1'b1;

  // instantiate function_92 for neuron804_1
  function_92 neuron804_1 (
      .a(input_layer[777]),
      .b(~input_layer[306]),
      .c(input_layer[1430]),
      .d(input_layer[824]),
      .e(input_layer[219]),
      .f(~input_layer[928]),
      .y(Y[804]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_274 for neuron805_1
  function_274 neuron805_1 (
      .a(input_layer[1373]),
      .b(~input_layer[1437]),
      .c(input_layer[1325]),
      .d(~input_layer[683]),
      .e(input_layer[1385]),
      .f(input_layer[640]),
      .y(Y[805]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_275 for neuron806_1
  function_275 neuron806_1 (
      .a(input_layer[145]),
      .b(input_layer[1098]),
      .c(input_layer[1392]),
      .d(input_layer[1500]),
      .e(~input_layer[730]),
      .f(~input_layer[1417]),
      .y(Y[806]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron807_1
  function_241 neuron807_1 (
      .a(input_layer[1430]),
      .b(~input_layer[747]),
      .c(input_layer[565]),
      .d(input_layer[513]),
      .e(input_layer[355]),
      .f(input_layer[293]),
      .y(Y[807]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron808_1
  function_67 neuron808_1 (
      .a(~input_layer[203]),
      .b(~input_layer[380]),
      .c(~input_layer[346]),
      .d(~input_layer[153]),
      .e(~input_layer[1157]),
      .y(Y[808]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_161 for neuron809_1
  function_161 neuron809_1 (
      .a(~input_layer[705]),
      .b(input_layer[482]),
      .c(~input_layer[634]),
      .d(~input_layer[352]),
      .e(input_layer[339]),
      .f(~input_layer[1403]),
      .y(Y[809]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_276 for neuron810_1
  function_276 neuron810_1 (
      .a(input_layer[260]),
      .b(~input_layer[506]),
      .c(input_layer[304]),
      .d(input_layer[688]),
      .e(input_layer[416]),
      .f(~input_layer[615]),
      .y(Y[810]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron811_1
  function_36 neuron811_1 (
      .a(input_layer[627]),
      .b(input_layer[548]),
      .c(input_layer[321]),
      .d(input_layer[124]),
      .e(~input_layer[373]),
      .f(input_layer[176]),
      .y(Y[811]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron812_1
  function_47 neuron812_1 (
      .a(input_layer[1494]),
      .b(input_layer[1243]),
      .c(input_layer[665]),
      .d(input_layer[90]),
      .e(input_layer[997]),
      .y(Y[812]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[813] = 1'b0;

  // instantiate function_124 for neuron814_1
  function_124 neuron814_1 (
      .a(~input_layer[1417]),
      .b(~input_layer[763]),
      .c(~input_layer[1436]),
      .d(~input_layer[1154]),
      .e(input_layer[532]),
      .f(~input_layer[798]),
      .y(Y[814]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron815_1
  function_84 neuron815_1 (
      .a(~input_layer[927]),
      .b(input_layer[1196]),
      .c(input_layer[1137]),
      .d(~input_layer[558]),
      .e(~input_layer[1557]),
      .y(Y[815]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron816_1
  function_39 neuron816_1 (
      .a(~input_layer[496]),
      .b(input_layer[1127]),
      .c(input_layer[1017]),
      .y(Y[816]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron817_1
  function_95 neuron817_1 (
      .a(input_layer[1420]),
      .b(~input_layer[1163]),
      .c(~input_layer[885]),
      .d(input_layer[210]),
      .y(Y[817]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron818_1
  function_1 neuron818_1 (
      .a(~input_layer[1428]),
      .b(~input_layer[1543]),
      .c(input_layer[861]),
      .d(input_layer[352]),
      .y(Y[818]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_277 for neuron819_1
  function_277 neuron819_1 (
      .a(input_layer[548]),
      .b(~input_layer[1237]),
      .c(~input_layer[73]),
      .d(~input_layer[99]),
      .e(input_layer[503]),
      .f(~input_layer[1406]),
      .y(Y[819]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron820_1
  function_27 neuron820_1 (
      .a(~input_layer[936]),
      .b(~input_layer[990]),
      .c(~input_layer[1295]),
      .y(Y[820]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron821_1
  function_27 neuron821_1 (
      .a(~input_layer[134]),
      .b(input_layer[753]),
      .c(~input_layer[1116]),
      .y(Y[821]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron822_1
  function_67 neuron822_1 (
      .a(~input_layer[183]),
      .b(~input_layer[564]),
      .c(~input_layer[257]),
      .d(input_layer[641]),
      .e(~input_layer[837]),
      .y(Y[822]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_278 for neuron823_1
  function_278 neuron823_1 (
      .a(~input_layer[1047]),
      .b(input_layer[491]),
      .c(input_layer[723]),
      .d(input_layer[645]),
      .e(~input_layer[1245]),
      .y(Y[823]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_279 for neuron824_1
  function_279 neuron824_1 (
      .a(input_layer[458]),
      .b(~input_layer[1082]),
      .c(~input_layer[1102]),
      .d(~input_layer[1090]),
      .e(input_layer[408]),
      .y(Y[824]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_124 for neuron825_1
  function_124 neuron825_1 (
      .a(~input_layer[1039]),
      .b(~input_layer[544]),
      .c(~input_layer[1023]),
      .d(input_layer[631]),
      .e(~input_layer[96]),
      .f(input_layer[698]),
      .y(Y[825]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron826_1
  function_63 neuron826_1 (
      .a(input_layer[1156]),
      .b(input_layer[512]),
      .c(~input_layer[318]),
      .d(~input_layer[535]),
      .e(input_layer[1084]),
      .y(Y[826]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_280 for neuron827_1
  function_280 neuron827_1 (
      .a(input_layer[199]),
      .b(~input_layer[360]),
      .c(input_layer[798]),
      .d(~input_layer[494]),
      .e(~input_layer[469]),
      .f(input_layer[261]),
      .y(Y[827]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_281 for neuron828_1
  function_281 neuron828_1 (
      .a(~input_layer[1131]),
      .b(~input_layer[1281]),
      .c(input_layer[697]),
      .d(input_layer[192]),
      .e(~input_layer[892]),
      .f(input_layer[618]),
      .y(Y[828]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron829_1
  function_17 neuron829_1 (
      .a(input_layer[1056]),
      .b(input_layer[500]),
      .c(input_layer[290]),
      .y(Y[829]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron830_1
  function_24 neuron830_1 (
      .a(~input_layer[1162]),
      .b(~input_layer[893]),
      .c(input_layer[217]),
      .y(Y[830]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron831_1
  function_67 neuron831_1 (
      .a(~input_layer[1416]),
      .b(input_layer[196]),
      .c(~input_layer[367]),
      .d(~input_layer[381]),
      .e(~input_layer[1474]),
      .y(Y[831]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron832_1
  function_36 neuron832_1 (
      .a(input_layer[890]),
      .b(input_layer[208]),
      .c(input_layer[1196]),
      .d(input_layer[375]),
      .e(input_layer[1254]),
      .f(input_layer[223]),
      .y(Y[832]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron833_1
  function_28 neuron833_1 (
      .a(~input_layer[406]),
      .b(~input_layer[236]),
      .c(~input_layer[201]),
      .d(~input_layer[1487]),
      .e(~input_layer[836]),
      .f(input_layer[1255]),
      .y(Y[833]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_282 for neuron834_1
  function_282 neuron834_1 (
      .a(input_layer[1030]),
      .b(~input_layer[1101]),
      .c(~input_layer[640]),
      .d(~input_layer[1305]),
      .e(~input_layer[863]),
      .f(input_layer[308]),
      .y(Y[834]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_269 for neuron835_1
  function_269 neuron835_1 (
      .a(input_layer[1540]),
      .b(~input_layer[833]),
      .c(input_layer[87]),
      .d(~input_layer[688]),
      .e(input_layer[1406]),
      .f(input_layer[1109]),
      .y(Y[835]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron836_1
  function_3 neuron836_1 (
      .a(~input_layer[974]),
      .b(~input_layer[751]),
      .c(~input_layer[1528]),
      .d(~input_layer[696]),
      .y(Y[836]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_283 for neuron837_1
  function_283 neuron837_1 (
      .a(input_layer[1171]),
      .b(input_layer[1042]),
      .c(~input_layer[664]),
      .d(~input_layer[277]),
      .e(~input_layer[614]),
      .f(~input_layer[670]),
      .y(Y[837]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_259 for neuron838_1
  function_259 neuron838_1 (
      .a(~input_layer[744]),
      .b(input_layer[1112]),
      .c(input_layer[1126]),
      .d(~input_layer[669]),
      .e(~input_layer[95]),
      .y(Y[838]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_275 for neuron839_1
  function_275 neuron839_1 (
      .a(~input_layer[538]),
      .b(input_layer[1271]),
      .c(input_layer[1273]),
      .d(input_layer[495]),
      .e(input_layer[1014]),
      .f(input_layer[1328]),
      .y(Y[839]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron840_1
  function_72 neuron840_1 (
      .a(input_layer[1221]),
      .b(~input_layer[1499]),
      .c(~input_layer[941]),
      .d(~input_layer[72]),
      .e(input_layer[1052]),
      .y(Y[840]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron841_1
  function_17 neuron841_1 (
      .a(input_layer[855]),
      .b(input_layer[240]),
      .c(input_layer[241]),
      .y(Y[841]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron842_1
  function_24 neuron842_1 (
      .a(~input_layer[308]),
      .b(~input_layer[991]),
      .c(~input_layer[870]),
      .y(Y[842]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_284 for neuron843_1
  function_284 neuron843_1 (
      .a(input_layer[487]),
      .b(~input_layer[256]),
      .c(input_layer[1478]),
      .d(input_layer[476]),
      .e(~input_layer[195]),
      .f(input_layer[787]),
      .y(Y[843]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron844_1
  function_27 neuron844_1 (
      .a(~input_layer[354]),
      .b(~input_layer[990]),
      .c(~input_layer[803]),
      .y(Y[844]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron845_1
  function_167 neuron845_1 (
      .a(input_layer[887]),
      .b(input_layer[1180]),
      .c(input_layer[1497]),
      .d(~input_layer[331]),
      .e(input_layer[259]),
      .y(Y[845]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron846_1
  function_26 neuron846_1 (
      .a(input_layer[1133]),
      .y(Y[846]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron847_1
  function_12 neuron847_1 (
      .a(~input_layer[253]),
      .b(input_layer[501]),
      .c(input_layer[98]),
      .y(Y[847]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_285 for neuron848_1
  function_285 neuron848_1 (
      .a(~input_layer[1479]),
      .b(input_layer[857]),
      .c(~input_layer[576]),
      .d(~input_layer[491]),
      .e(~input_layer[73]),
      .f(~input_layer[125]),
      .y(Y[848]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron849_1
  function_286 neuron849_1 (
      .a(input_layer[1183]),
      .b(~input_layer[620]),
      .c(input_layer[1351]),
      .d(~input_layer[121]),
      .e(~input_layer[69]),
      .y(Y[849]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_287 for neuron850_1
  function_287 neuron850_1 (
      .a(~input_layer[544]),
      .b(input_layer[329]),
      .c(input_layer[1367]),
      .d(input_layer[1244]),
      .e(~input_layer[562]),
      .f(~input_layer[794]),
      .y(Y[850]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron851_1
  function_52 neuron851_1 (
      .a(input_layer[250]),
      .b(~input_layer[695]),
      .c(~input_layer[825]),
      .d(~input_layer[1555]),
      .e(input_layer[66]),
      .f(~input_layer[281]),
      .y(Y[851]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron852_1
  function_149 neuron852_1 (
      .a(~input_layer[1486]),
      .b(input_layer[365]),
      .c(input_layer[1058]),
      .d(~input_layer[548]),
      .y(Y[852]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron853_1
  function_28 neuron853_1 (
      .a(~input_layer[582]),
      .b(~input_layer[1018]),
      .c(~input_layer[1486]),
      .d(~input_layer[1476]),
      .e(~input_layer[1332]),
      .f(~input_layer[946]),
      .y(Y[853]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron854_1
  function_62 neuron854_1 (
      .a(input_layer[1167]),
      .b(~input_layer[651]),
      .c(input_layer[1324]),
      .d(input_layer[290]),
      .e(input_layer[1293]),
      .f(~input_layer[520]),
      .y(Y[854]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron855_1
  function_214 neuron855_1 (
      .a(input_layer[192]),
      .b(input_layer[566]),
      .c(~input_layer[474]),
      .d(input_layer[451]),
      .e(input_layer[1141]),
      .f(input_layer[163]),
      .y(Y[855]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron856_1
  function_167 neuron856_1 (
      .a(~input_layer[645]),
      .b(input_layer[1477]),
      .c(input_layer[1420]),
      .d(input_layer[513]),
      .e(input_layer[158]),
      .y(Y[856]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[857] = 1'b1;

  // instantiate function_24 for neuron858_1
  function_24 neuron858_1 (
      .a(~input_layer[639]),
      .b(~input_layer[578]),
      .c(input_layer[1447]),
      .y(Y[858]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_247 for neuron859_1
  function_247 neuron859_1 (
      .a(input_layer[1227]),
      .b(input_layer[856]),
      .c(input_layer[233]),
      .d(~input_layer[712]),
      .e(input_layer[1277]),
      .f(~input_layer[382]),
      .y(Y[859]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron860_1
  function_113 neuron860_1 (
      .a(input_layer[1152]),
      .b(input_layer[826]),
      .c(~input_layer[633]),
      .d(input_layer[396]),
      .e(input_layer[619]),
      .y(Y[860]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_288 for neuron861_1
  function_288 neuron861_1 (
      .a(~input_layer[692]),
      .b(input_layer[1113]),
      .c(~input_layer[214]),
      .d(~input_layer[1237]),
      .e(input_layer[536]),
      .f(input_layer[1244]),
      .y(Y[861]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron862_1
  function_27 neuron862_1 (
      .a(~input_layer[255]),
      .b(~input_layer[1079]),
      .c(~input_layer[883]),
      .y(Y[862]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_289 for neuron863_1
  function_289 neuron863_1 (
      .a(~input_layer[1413]),
      .b(~input_layer[564]),
      .c(input_layer[521]),
      .d(~input_layer[934]),
      .e(~input_layer[823]),
      .f(input_layer[714]),
      .y(Y[863]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron864_1
  function_3 neuron864_1 (
      .a(~input_layer[460]),
      .b(~input_layer[946]),
      .c(~input_layer[1268]),
      .d(~input_layer[1542]),
      .y(Y[864]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron865_1
  function_290 neuron865_1 (
      .a(~input_layer[932]),
      .b(~input_layer[546]),
      .c(input_layer[307]),
      .d(~input_layer[422]),
      .e(~input_layer[478]),
      .f(~input_layer[1092]),
      .y(Y[865]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_291 for neuron866_1
  function_291 neuron866_1 (
      .a(input_layer[1225]),
      .b(~input_layer[128]),
      .c(~input_layer[83]),
      .d(input_layer[1022]),
      .e(input_layer[1552]),
      .y(Y[866]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron867_1
  function_17 neuron867_1 (
      .a(input_layer[914]),
      .b(input_layer[819]),
      .c(input_layer[859]),
      .y(Y[867]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron868_1
  function_35 neuron868_1 (
      .a(~input_layer[582]),
      .b(~input_layer[1070]),
      .c(input_layer[811]),
      .d(~input_layer[158]),
      .e(input_layer[1035]),
      .y(Y[868]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron869_1
  function_119 neuron869_1 (
      .a(~input_layer[1137]),
      .b(~input_layer[1102]),
      .c(~input_layer[825]),
      .d(input_layer[589]),
      .e(~input_layer[374]),
      .y(Y[869]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron870_1
  function_47 neuron870_1 (
      .a(input_layer[1048]),
      .b(input_layer[796]),
      .c(input_layer[775]),
      .d(~input_layer[811]),
      .e(input_layer[1052]),
      .y(Y[870]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron871_1
  function_0 neuron871_1 (
      .a(~input_layer[510]),
      .b(~input_layer[665]),
      .c(~input_layer[1352]),
      .d(input_layer[667]),
      .e(input_layer[275]),
      .y(Y[871]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron872_1
  function_8 neuron872_1 (
      .a(input_layer[976]),
      .b(input_layer[511]),
      .c(input_layer[925]),
      .d(~input_layer[424]),
      .y(Y[872]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_292 for neuron873_1
  function_292 neuron873_1 (
      .a(~input_layer[638]),
      .b(~input_layer[1050]),
      .c(~input_layer[95]),
      .d(input_layer[1041]),
      .e(input_layer[1502]),
      .f(input_layer[1284]),
      .y(Y[873]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[874] = 1'b0;

  // instantiate function_235 for neuron875_1
  function_235 neuron875_1 (
      .a(~input_layer[706]),
      .b(~input_layer[1282]),
      .c(~input_layer[140]),
      .d(~input_layer[1163]),
      .e(input_layer[1558]),
      .y(Y[875]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron876_1
  function_29 neuron876_1 (
      .a(~input_layer[870]),
      .b(~input_layer[1439]),
      .y(Y[876]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron877_1
  function_29 neuron877_1 (
      .a(~input_layer[1162]),
      .b(~input_layer[569]),
      .y(Y[877]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_166 for neuron878_1
  function_166 neuron878_1 (
      .a(input_layer[1277]),
      .b(~input_layer[860]),
      .c(~input_layer[210]),
      .d(~input_layer[85]),
      .e(~input_layer[438]),
      .f(~input_layer[1042]),
      .y(Y[878]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_173 for neuron879_1
  function_173 neuron879_1 (
      .a(~input_layer[316]),
      .b(input_layer[1274]),
      .c(~input_layer[1545]),
      .d(~input_layer[514]),
      .e(~input_layer[1091]),
      .y(Y[879]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_293 for neuron880_1
  function_293 neuron880_1 (
      .a(~input_layer[634]),
      .b(~input_layer[153]),
      .c(input_layer[535]),
      .d(input_layer[563]),
      .e(input_layer[1522]),
      .f(~input_layer[1449]),
      .y(Y[880]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron881_1
  function_21 neuron881_1 (
      .a(input_layer[371]),
      .b(input_layer[295]),
      .c(~input_layer[1423]),
      .d(~input_layer[1321]),
      .e(~input_layer[478]),
      .y(Y[881]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron882_1
  function_57 neuron882_1 (
      .a(input_layer[1142]),
      .b(input_layer[1359]),
      .c(~input_layer[1178]),
      .d(~input_layer[101]),
      .e(~input_layer[571]),
      .f(~input_layer[226]),
      .y(Y[882]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron883_1
  function_55 neuron883_1 (
      .a(~input_layer[687]),
      .b(~input_layer[740]),
      .c(~input_layer[880]),
      .d(input_layer[293]),
      .e(input_layer[1213]),
      .y(Y[883]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron884_1
  function_57 neuron884_1 (
      .a(~input_layer[818]),
      .b(input_layer[589]),
      .c(~input_layer[1357]),
      .d(~input_layer[508]),
      .e(input_layer[575]),
      .f(input_layer[102]),
      .y(Y[884]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_294 for neuron885_1
  function_294 neuron885_1 (
      .a(input_layer[554]),
      .b(~input_layer[650]),
      .c(~input_layer[382]),
      .d(input_layer[702]),
      .e(input_layer[960]),
      .f(~input_layer[823]),
      .y(Y[885]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron886_1
  function_36 neuron886_1 (
      .a(input_layer[947]),
      .b(input_layer[1329]),
      .c(input_layer[363]),
      .d(input_layer[690]),
      .e(input_layer[122]),
      .f(~input_layer[1521]),
      .y(Y[886]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron887_1
  function_167 neuron887_1 (
      .a(input_layer[185]),
      .b(input_layer[1198]),
      .c(~input_layer[908]),
      .d(~input_layer[930]),
      .e(~input_layer[916]),
      .y(Y[887]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron888_1
  function_3 neuron888_1 (
      .a(~input_layer[1420]),
      .b(~input_layer[935]),
      .c(~input_layer[546]),
      .d(input_layer[419]),
      .y(Y[888]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron889_1
  function_48 neuron889_1 (
      .a(input_layer[1189]),
      .b(input_layer[304]),
      .c(input_layer[864]),
      .d(input_layer[84]),
      .e(input_layer[497]),
      .y(Y[889]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron890_1
  function_39 neuron890_1 (
      .a(~input_layer[1142]),
      .b(input_layer[1420]),
      .c(~input_layer[1004]),
      .y(Y[890]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_103 for neuron891_1
  function_103 neuron891_1 (
      .a(input_layer[1323]),
      .b(~input_layer[203]),
      .c(input_layer[700]),
      .d(input_layer[1324]),
      .e(input_layer[1125]),
      .f(~input_layer[1006]),
      .y(Y[891]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron892_1
  function_30 neuron892_1 (
      .a(input_layer[765]),
      .b(~input_layer[607]),
      .c(input_layer[217]),
      .d(input_layer[355]),
      .y(Y[892]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_295 for neuron893_1
  function_295 neuron893_1 (
      .a(input_layer[439]),
      .b(~input_layer[816]),
      .c(~input_layer[1445]),
      .d(~input_layer[353]),
      .e(~input_layer[931]),
      .f(~input_layer[891]),
      .y(Y[893]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron894_1
  function_16 neuron894_1 (
      .a(input_layer[749]),
      .b(input_layer[1136]),
      .y(Y[894]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron895_1
  function_128 neuron895_1 (
      .a(~input_layer[864]),
      .b(input_layer[621]),
      .c(~input_layer[445]),
      .d(~input_layer[1248]),
      .y(Y[895]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron896_1
  function_30 neuron896_1 (
      .a(input_layer[468]),
      .b(input_layer[1386]),
      .c(input_layer[1316]),
      .d(input_layer[333]),
      .y(Y[896]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron897_1
  function_39 neuron897_1 (
      .a(~input_layer[1482]),
      .b(input_layer[1031]),
      .c(input_layer[1275]),
      .y(Y[897]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron898_1
  function_3 neuron898_1 (
      .a(~input_layer[517]),
      .b(~input_layer[746]),
      .c(~input_layer[1052]),
      .d(~input_layer[798]),
      .y(Y[898]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_296 for neuron899_1
  function_296 neuron899_1 (
      .a(input_layer[704]),
      .b(input_layer[874]),
      .c(input_layer[1389]),
      .d(~input_layer[1524]),
      .e(input_layer[571]),
      .f(~input_layer[411]),
      .y(Y[899]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron900_1
  function_126 neuron900_1 (
      .a(~input_layer[191]),
      .b(~input_layer[1137]),
      .c(~input_layer[912]),
      .d(input_layer[534]),
      .e(~input_layer[94]),
      .y(Y[900]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron901_1
  function_27 neuron901_1 (
      .a(~input_layer[1111]),
      .b(~input_layer[545]),
      .c(~input_layer[544]),
      .y(Y[901]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron902_1
  function_25 neuron902_1 (
      .a(input_layer[185]),
      .b(input_layer[1491]),
      .c(~input_layer[719]),
      .d(input_layer[387]),
      .e(input_layer[413]),
      .y(Y[902]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron903_1
  function_27 neuron903_1 (
      .a(~input_layer[1089]),
      .b(~input_layer[1093]),
      .c(~input_layer[600]),
      .y(Y[903]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron904_1
  function_4 neuron904_1 (
      .a(input_layer[538]),
      .b(~input_layer[1169]),
      .c(~input_layer[994]),
      .d(~input_layer[848]),
      .e(~input_layer[901]),
      .y(Y[904]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_297 for neuron905_1
  function_297 neuron905_1 (
      .a(~input_layer[1242]),
      .b(input_layer[1495]),
      .c(~input_layer[214]),
      .d(input_layer[76]),
      .e(~input_layer[151]),
      .f(~input_layer[138]),
      .y(Y[905]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_211 for neuron906_1
  function_211 neuron906_1 (
      .a(~input_layer[440]),
      .b(~input_layer[798]),
      .c(input_layer[1170]),
      .d(input_layer[252]),
      .e(~input_layer[1311]),
      .f(~input_layer[536]),
      .y(Y[906]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron907_1
  function_60 neuron907_1 (
      .a(input_layer[1113]),
      .b(~input_layer[350]),
      .c(~input_layer[1408]),
      .d(~input_layer[358]),
      .e(input_layer[1199]),
      .y(Y[907]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron908_1
  function_19 neuron908_1 (
      .a(~input_layer[418]),
      .b(~input_layer[130]),
      .c(~input_layer[1099]),
      .d(input_layer[1069]),
      .y(Y[908]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron909_1
  function_17 neuron909_1 (
      .a(input_layer[142]),
      .b(input_layer[1313]),
      .c(input_layer[1544]),
      .y(Y[909]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron910_1
  function_119 neuron910_1 (
      .a(~input_layer[320]),
      .b(input_layer[474]),
      .c(input_layer[1336]),
      .d(input_layer[14]),
      .e(~input_layer[1010]),
      .y(Y[910]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron911_1
  function_107 neuron911_1 (
      .a(~input_layer[609]),
      .b(~input_layer[947]),
      .c(input_layer[453]),
      .d(input_layer[1354]),
      .e(~input_layer[1413]),
      .y(Y[911]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_102 for neuron912_1
  function_102 neuron912_1 (
      .a(~input_layer[586]),
      .b(~input_layer[575]),
      .c(input_layer[482]),
      .d(input_layer[1192]),
      .e(~input_layer[451]),
      .f(~input_layer[853]),
      .y(Y[912]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron913_1
  function_298 neuron913_1 (
      .a(~input_layer[513]),
      .b(input_layer[501]),
      .c(~input_layer[1172]),
      .d(~input_layer[1224]),
      .e(~input_layer[360]),
      .f(~input_layer[1009]),
      .y(Y[913]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron914_1
  function_49 neuron914_1 (
      .a(input_layer[252]),
      .b(~input_layer[1418]),
      .c(input_layer[1087]),
      .d(~input_layer[1534]),
      .e(~input_layer[1549]),
      .y(Y[914]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron915_1
  function_165 neuron915_1 (
      .a(~input_layer[200]),
      .b(input_layer[497]),
      .c(~input_layer[180]),
      .d(input_layer[704]),
      .e(input_layer[1260]),
      .y(Y[915]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron916_1
  function_8 neuron916_1 (
      .a(input_layer[1076]),
      .b(input_layer[1222]),
      .c(input_layer[239]),
      .d(~input_layer[1148]),
      .y(Y[916]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_273 for neuron917_1
  function_273 neuron917_1 (
      .a(input_layer[831]),
      .b(~input_layer[1189]),
      .c(~input_layer[1500]),
      .d(~input_layer[483]),
      .e(~input_layer[484]),
      .y(Y[917]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron918_1
  function_95 neuron918_1 (
      .a(input_layer[1487]),
      .b(~input_layer[1155]),
      .c(input_layer[520]),
      .d(~input_layer[1352]),
      .y(Y[918]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron919_1
  function_36 neuron919_1 (
      .a(input_layer[462]),
      .b(input_layer[445]),
      .c(~input_layer[922]),
      .d(input_layer[371]),
      .e(input_layer[906]),
      .f(input_layer[154]),
      .y(Y[919]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[920] = 1'b0;

  // instantiate function_214 for neuron921_1
  function_214 neuron921_1 (
      .a(input_layer[1430]),
      .b(input_layer[885]),
      .c(input_layer[1489]),
      .d(input_layer[1375]),
      .e(input_layer[1522]),
      .f(~input_layer[1007]),
      .y(Y[921]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron922_1
  function_248 neuron922_1 (
      .a(input_layer[927]),
      .b(~input_layer[509]),
      .c(input_layer[403]),
      .d(~input_layer[370]),
      .e(~input_layer[502]),
      .f(~input_layer[217]),
      .y(Y[922]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron923_1
  function_299 neuron923_1 (
      .a(~input_layer[1208]),
      .b(~input_layer[88]),
      .c(input_layer[931]),
      .d(~input_layer[822]),
      .e(~input_layer[249]),
      .y(Y[923]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_50 for neuron924_1
  function_50 neuron924_1 (
      .a(input_layer[747]),
      .b(input_layer[621]),
      .c(~input_layer[1252]),
      .d(~input_layer[321]),
      .e(input_layer[784]),
      .f(input_layer[393]),
      .y(Y[924]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_300 for neuron925_1
  function_300 neuron925_1 (
      .a(~input_layer[752]),
      .b(input_layer[475]),
      .c(input_layer[1142]),
      .d(input_layer[1192]),
      .e(~input_layer[306]),
      .y(Y[925]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron926_1
  function_67 neuron926_1 (
      .a(~input_layer[187]),
      .b(~input_layer[1088]),
      .c(input_layer[582]),
      .d(input_layer[1524]),
      .e(~input_layer[604]),
      .y(Y[926]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[927] = 1'b1;

  // instantiate function_167 for neuron928_1
  function_167 neuron928_1 (
      .a(input_layer[252]),
      .b(input_layer[1254]),
      .c(input_layer[208]),
      .d(~input_layer[826]),
      .e(input_layer[528]),
      .y(Y[928]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron929_1
  function_26 neuron929_1 (
      .a(input_layer[636]),
      .y(Y[929]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron930_1
  function_112 neuron930_1 (
      .a(input_layer[719]),
      .b(~input_layer[793]),
      .c(input_layer[691]),
      .d(~input_layer[557]),
      .e(~input_layer[494]),
      .f(input_layer[247]),
      .y(Y[930]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron931_1
  function_121 neuron931_1 (
      .a(~input_layer[486]),
      .b(input_layer[151]),
      .c(input_layer[88]),
      .d(input_layer[809]),
      .e(~input_layer[1020]),
      .y(Y[931]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron932_1
  function_27 neuron932_1 (
      .a(~input_layer[298]),
      .b(~input_layer[310]),
      .c(input_layer[982]),
      .y(Y[932]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron933_1
  function_33 neuron933_1 (
      .a(~input_layer[987]),
      .b(~input_layer[470]),
      .c(input_layer[1293]),
      .d(input_layer[587]),
      .e(input_layer[920]),
      .f(~input_layer[45]),
      .y(Y[933]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_301 for neuron934_1
  function_301 neuron934_1 (
      .a(input_layer[742]),
      .b(~input_layer[1260]),
      .c(input_layer[316]),
      .d(~input_layer[1257]),
      .e(~input_layer[166]),
      .f(input_layer[284]),
      .y(Y[934]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron935_1
  function_46 neuron935_1 (
      .a(input_layer[922]),
      .b(input_layer[363]),
      .c(input_layer[261]),
      .d(~input_layer[1489]),
      .e(input_layer[1265]),
      .y(Y[935]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron936_1
  function_70 neuron936_1 (
      .a(~input_layer[1417]),
      .b(~input_layer[1482]),
      .c(~input_layer[77]),
      .d(~input_layer[1503]),
      .e(~input_layer[467]),
      .f(input_layer[13]),
      .y(Y[936]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron937_1
  function_46 neuron937_1 (
      .a(input_layer[1317]),
      .b(input_layer[349]),
      .c(~input_layer[272]),
      .d(input_layer[585]),
      .e(input_layer[285]),
      .y(Y[937]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron938_1
  function_8 neuron938_1 (
      .a(input_layer[811]),
      .b(input_layer[959]),
      .c(input_layer[77]),
      .d(~input_layer[1245]),
      .y(Y[938]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron939_1
  function_95 neuron939_1 (
      .a(~input_layer[1191]),
      .b(input_layer[1310]),
      .c(input_layer[1013]),
      .d(~input_layer[178]),
      .y(Y[939]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron940_1
  function_55 neuron940_1 (
      .a(~input_layer[553]),
      .b(~input_layer[1470]),
      .c(~input_layer[1548]),
      .d(input_layer[300]),
      .e(~input_layer[1529]),
      .y(Y[940]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron941_1
  function_84 neuron941_1 (
      .a(~input_layer[592]),
      .b(~input_layer[661]),
      .c(input_layer[134]),
      .d(~input_layer[773]),
      .e(input_layer[298]),
      .y(Y[941]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_98 for neuron942_1
  function_98 neuron942_1 (
      .a(~input_layer[793]),
      .b(~input_layer[937]),
      .c(~input_layer[873]),
      .d(~input_layer[695]),
      .e(input_layer[1028]),
      .f(~input_layer[188]),
      .y(Y[942]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron943_1
  function_29 neuron943_1 (
      .a(~input_layer[1133]),
      .b(~input_layer[1180]),
      .y(Y[943]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron944_1
  function_12 neuron944_1 (
      .a(input_layer[1074]),
      .b(~input_layer[319]),
      .c(input_layer[299]),
      .y(Y[944]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron945_1
  function_6 neuron945_1 (
      .a(~input_layer[327]),
      .b(input_layer[428]),
      .c(input_layer[1429]),
      .d(input_layer[837]),
      .e(input_layer[1002]),
      .f(input_layer[115]),
      .y(Y[945]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron946_1
  function_39 neuron946_1 (
      .a(input_layer[238]),
      .b(~input_layer[657]),
      .c(input_layer[647]),
      .y(Y[946]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_302 for neuron947_1
  function_302 neuron947_1 (
      .a(input_layer[496]),
      .b(~input_layer[975]),
      .c(~input_layer[301]),
      .d(input_layer[481]),
      .e(~input_layer[306]),
      .f(~input_layer[993]),
      .y(Y[947]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron948_1
  function_90 neuron948_1 (
      .a(~input_layer[852]),
      .b(~input_layer[1153]),
      .c(input_layer[633]),
      .d(~input_layer[1042]),
      .e(~input_layer[1552]),
      .y(Y[948]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_236 for neuron949_1
  function_236 neuron949_1 (
      .a(input_layer[917]),
      .b(input_layer[723]),
      .c(input_layer[976]),
      .d(input_layer[861]),
      .e(input_layer[260]),
      .f(~input_layer[844]),
      .y(Y[949]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron950_1
  function_67 neuron950_1 (
      .a(~input_layer[1107]),
      .b(~input_layer[403]),
      .c(~input_layer[1474]),
      .d(~input_layer[196]),
      .e(~input_layer[493]),
      .y(Y[950]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_164 for neuron951_1
  function_164 neuron951_1 (
      .a(~input_layer[1186]),
      .b(~input_layer[1192]),
      .c(~input_layer[1078]),
      .d(~input_layer[605]),
      .e(~input_layer[1090]),
      .f(~input_layer[283]),
      .y(Y[951]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron952_1
  function_24 neuron952_1 (
      .a(~input_layer[1083]),
      .b(input_layer[748]),
      .c(input_layer[862]),
      .y(Y[952]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron953_1
  function_36 neuron953_1 (
      .a(input_layer[310]),
      .b(input_layer[378]),
      .c(input_layer[621]),
      .d(input_layer[1224]),
      .e(input_layer[1269]),
      .f(input_layer[1553]),
      .y(Y[953]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron954_1
  function_299 neuron954_1 (
      .a(~input_layer[555]),
      .b(input_layer[607]),
      .c(~input_layer[651]),
      .d(input_layer[608]),
      .e(~input_layer[1543]),
      .y(Y[954]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron955_1
  function_78 neuron955_1 (
      .a(~input_layer[630]),
      .b(~input_layer[1002]),
      .c(~input_layer[262]),
      .d(input_layer[1259]),
      .e(~input_layer[1021]),
      .f(~input_layer[27]),
      .y(Y[955]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron956_1
  function_42 neuron956_1 (
      .a(input_layer[1369]),
      .b(input_layer[1300]),
      .c(~input_layer[978]),
      .d(input_layer[566]),
      .y(Y[956]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron957_1
  function_27 neuron957_1 (
      .a(~input_layer[327]),
      .b(~input_layer[1496]),
      .c(~input_layer[949]),
      .y(Y[957]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron958_1
  function_26 neuron958_1 (
      .a(~input_layer[874]),
      .y(Y[958]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron959_1
  function_155 neuron959_1 (
      .a(~input_layer[1046]),
      .b(~input_layer[1313]),
      .c(~input_layer[1072]),
      .d(~input_layer[195]),
      .e(~input_layer[569]),
      .f(~input_layer[1281]),
      .y(Y[959]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron960_1
  function_3 neuron960_1 (
      .a(~input_layer[365]),
      .b(~input_layer[1528]),
      .c(~input_layer[498]),
      .d(~input_layer[363]),
      .y(Y[960]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron961_1
  function_186 neuron961_1 (
      .a(~input_layer[1031]),
      .b(input_layer[943]),
      .c(~input_layer[611]),
      .d(~input_layer[356]),
      .y(Y[961]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron962_1
  function_303 neuron962_1 (
      .a(input_layer[816]),
      .b(input_layer[1432]),
      .c(~input_layer[999]),
      .d(input_layer[506]),
      .e(~input_layer[261]),
      .f(input_layer[1557]),
      .y(Y[962]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron963_1
  function_24 neuron963_1 (
      .a(~input_layer[854]),
      .b(~input_layer[849]),
      .c(input_layer[297]),
      .y(Y[963]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_304 for neuron964_1
  function_304 neuron964_1 (
      .a(~input_layer[865]),
      .b(input_layer[544]),
      .c(input_layer[551]),
      .d(~input_layer[893]),
      .e(~input_layer[1052]),
      .f(input_layer[1148]),
      .y(Y[964]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron965_1
  function_14 neuron965_1 (
      .a(input_layer[153]),
      .b(~input_layer[482]),
      .c(~input_layer[400]),
      .d(input_layer[94]),
      .e(input_layer[853]),
      .f(input_layer[88]),
      .y(Y[965]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron966_1
  function_29 neuron966_1 (
      .a(~input_layer[720]),
      .b(~input_layer[566]),
      .y(Y[966]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron967_1
  function_29 neuron967_1 (
      .a(~input_layer[1111]),
      .b(~input_layer[1214]),
      .y(Y[967]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron968_1
  function_46 neuron968_1 (
      .a(input_layer[1243]),
      .b(input_layer[947]),
      .c(input_layer[779]),
      .d(~input_layer[1335]),
      .e(input_layer[670]),
      .y(Y[968]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron969_1
  function_36 neuron969_1 (
      .a(input_layer[714]),
      .b(input_layer[1410]),
      .c(input_layer[159]),
      .d(~input_layer[1196]),
      .e(input_layer[458]),
      .f(~input_layer[17]),
      .y(Y[969]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron970_1
  function_241 neuron970_1 (
      .a(input_layer[421]),
      .b(input_layer[1241]),
      .c(~input_layer[872]),
      .d(input_layer[181]),
      .e(input_layer[891]),
      .f(input_layer[733]),
      .y(Y[970]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron971_1
  function_8 neuron971_1 (
      .a(input_layer[143]),
      .b(~input_layer[912]),
      .c(input_layer[356]),
      .d(input_layer[351]),
      .y(Y[971]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[972] = 1'b0;

  // instantiate function_305 for neuron973_1
  function_305 neuron973_1 (
      .a(~input_layer[609]),
      .b(~input_layer[492]),
      .c(input_layer[1113]),
      .d(~input_layer[937]),
      .e(input_layer[1495]),
      .y(Y[973]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron974_1
  function_92 neuron974_1 (
      .a(input_layer[300]),
      .b(input_layer[1488]),
      .c(input_layer[1364]),
      .d(input_layer[837]),
      .e(~input_layer[1207]),
      .f(input_layer[1031]),
      .y(Y[974]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_127 for neuron975_1
  function_127 neuron975_1 (
      .a(input_layer[1091]),
      .b(input_layer[1222]),
      .c(input_layer[212]),
      .d(~input_layer[605]),
      .e(~input_layer[1103]),
      .f(~input_layer[1349]),
      .y(Y[975]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_306 for neuron976_1
  function_306 neuron976_1 (
      .a(~input_layer[708]),
      .b(~input_layer[1542]),
      .c(~input_layer[790]),
      .d(~input_layer[1479]),
      .e(input_layer[385]),
      .f(input_layer[1325]),
      .y(Y[976]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron977_1
  function_74 neuron977_1 (
      .a(input_layer[1089]),
      .b(~input_layer[720]),
      .c(~input_layer[657]),
      .d(input_layer[815]),
      .e(input_layer[1330]),
      .f(input_layer[537]),
      .y(Y[977]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron978_1
  function_48 neuron978_1 (
      .a(input_layer[149]),
      .b(input_layer[1190]),
      .c(input_layer[182]),
      .d(input_layer[1012]),
      .e(input_layer[334]),
      .y(Y[978]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron979_1
  function_307 neuron979_1 (
      .a(input_layer[312]),
      .b(input_layer[1018]),
      .c(~input_layer[567]),
      .d(~input_layer[1360]),
      .e(~input_layer[1259]),
      .y(Y[979]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron980_1
  function_179 neuron980_1 (
      .a(input_layer[327]),
      .b(~input_layer[1052]),
      .c(~input_layer[1087]),
      .d(~input_layer[1542]),
      .e(~input_layer[528]),
      .y(Y[980]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron981_1
  function_113 neuron981_1 (
      .a(~input_layer[760]),
      .b(~input_layer[1317]),
      .c(~input_layer[309]),
      .d(~input_layer[1254]),
      .e(input_layer[1445]),
      .y(Y[981]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron982_1
  function_126 neuron982_1 (
      .a(~input_layer[356]),
      .b(~input_layer[264]),
      .c(input_layer[459]),
      .d(~input_layer[833]),
      .e(~input_layer[93]),
      .y(Y[982]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron983_1
  function_17 neuron983_1 (
      .a(input_layer[1135]),
      .b(input_layer[642]),
      .c(input_layer[269]),
      .y(Y[983]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron984_1
  function_35 neuron984_1 (
      .a(~input_layer[130]),
      .b(~input_layer[1239]),
      .c(~input_layer[77]),
      .d(input_layer[406]),
      .e(input_layer[731]),
      .y(Y[984]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron985_1
  function_44 neuron985_1 (
      .a(~input_layer[1416]),
      .b(~input_layer[1152]),
      .c(input_layer[403]),
      .d(input_layer[243]),
      .e(input_layer[241]),
      .y(Y[985]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_308 for neuron986_1
  function_308 neuron986_1 (
      .a(~input_layer[152]),
      .b(input_layer[592]),
      .c(input_layer[409]),
      .d(~input_layer[887]),
      .e(~input_layer[1381]),
      .f(input_layer[932]),
      .y(Y[986]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron987_1
  function_35 neuron987_1 (
      .a(~input_layer[1490]),
      .b(input_layer[593]),
      .c(~input_layer[1282]),
      .d(input_layer[1305]),
      .e(~input_layer[1428]),
      .y(Y[987]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron988_1
  function_67 neuron988_1 (
      .a(~input_layer[192]),
      .b(~input_layer[991]),
      .c(~input_layer[188]),
      .d(~input_layer[1044]),
      .e(input_layer[802]),
      .y(Y[988]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron989_1
  function_67 neuron989_1 (
      .a(~input_layer[416]),
      .b(~input_layer[965]),
      .c(~input_layer[743]),
      .d(~input_layer[1095]),
      .e(~input_layer[1446]),
      .y(Y[989]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron990_1
  function_70 neuron990_1 (
      .a(~input_layer[203]),
      .b(~input_layer[1034]),
      .c(input_layer[623]),
      .d(~input_layer[1256]),
      .e(~input_layer[178]),
      .f(~input_layer[1459]),
      .y(Y[990]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_309 for neuron991_1
  function_309 neuron991_1 (
      .a(input_layer[441]),
      .b(~input_layer[132]),
      .c(~input_layer[976]),
      .d(~input_layer[742]),
      .e(input_layer[1197]),
      .f(~input_layer[318]),
      .y(Y[991]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron992_1
  function_26 neuron992_1 (
      .a(input_layer[920]),
      .y(Y[992]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_310 for neuron993_1
  function_310 neuron993_1 (
      .a(~input_layer[1055]),
      .b(~input_layer[389]),
      .c(input_layer[577]),
      .d(input_layer[685]),
      .e(~input_layer[1153]),
      .f(input_layer[786]),
      .y(Y[993]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_311 for neuron994_1
  function_311 neuron994_1 (
      .a(~input_layer[291]),
      .b(input_layer[1492]),
      .c(~input_layer[1265]),
      .d(~input_layer[1527]),
      .e(~input_layer[75]),
      .f(input_layer[791]),
      .y(Y[994]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron995_1
  function_183 neuron995_1 (
      .a(~input_layer[371]),
      .b(input_layer[720]),
      .c(input_layer[1209]),
      .d(~input_layer[957]),
      .e(input_layer[24]),
      .f(~input_layer[952]),
      .y(Y[995]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron996_1
  function_48 neuron996_1 (
      .a(input_layer[313]),
      .b(input_layer[79]),
      .c(input_layer[86]),
      .d(~input_layer[861]),
      .e(input_layer[838]),
      .y(Y[996]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_312 for neuron997_1
  function_312 neuron997_1 (
      .a(~input_layer[661]),
      .b(input_layer[404]),
      .c(input_layer[290]),
      .d(~input_layer[82]),
      .e(~input_layer[1173]),
      .f(~input_layer[1567]),
      .y(Y[997]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron998_1
  function_0 neuron998_1 (
      .a(~input_layer[1141]),
      .b(~input_layer[535]),
      .c(~input_layer[589]),
      .d(input_layer[866]),
      .e(~input_layer[702]),
      .y(Y[998]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_313 for neuron999_1
  function_313 neuron999_1 (
      .a(input_layer[908]),
      .b(~input_layer[1391]),
      .c(~input_layer[637]),
      .d(~input_layer[546]),
      .e(~input_layer[871]),
      .f(input_layer[103]),
      .y(Y[999]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_305 for neuron1000_1
  function_305 neuron1000_1 (
      .a(~input_layer[520]),
      .b(~input_layer[157]),
      .c(input_layer[443]),
      .d(~input_layer[97]),
      .e(input_layer[960]),
      .y(Y[1000]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1001_1
  function_172 neuron1001_1 (
      .a(~input_layer[1487]),
      .b(~input_layer[1419]),
      .c(~input_layer[1259]),
      .d(~input_layer[1001]),
      .e(~input_layer[1048]),
      .f(input_layer[432]),
      .y(Y[1001]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1002_1
  function_19 neuron1002_1 (
      .a(~input_layer[703]),
      .b(~input_layer[610]),
      .c(input_layer[416]),
      .d(~input_layer[300]),
      .y(Y[1002]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1003_1
  function_87 neuron1003_1 (
      .a(input_layer[716]),
      .b(input_layer[1422]),
      .c(~input_layer[944]),
      .d(~input_layer[350]),
      .e(~input_layer[451]),
      .y(Y[1003]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1004_1
  function_3 neuron1004_1 (
      .a(~input_layer[657]),
      .b(~input_layer[493]),
      .c(input_layer[925]),
      .d(~input_layer[1441]),
      .y(Y[1004]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron1005_1
  function_70 neuron1005_1 (
      .a(~input_layer[1316]),
      .b(~input_layer[1480]),
      .c(input_layer[837]),
      .d(~input_layer[397]),
      .e(input_layer[1101]),
      .f(~input_layer[1008]),
      .y(Y[1005]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_314 for neuron1006_1
  function_314 neuron1006_1 (
      .a(input_layer[542]),
      .b(~input_layer[754]),
      .c(input_layer[422]),
      .d(input_layer[586]),
      .e(~input_layer[217]),
      .y(Y[1006]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1007_1
  function_48 neuron1007_1 (
      .a(input_layer[913]),
      .b(input_layer[1483]),
      .c(input_layer[1496]),
      .d(input_layer[374]),
      .e(input_layer[1148]),
      .y(Y[1007]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron1008_1
  function_157 neuron1008_1 (
      .a(input_layer[760]),
      .b(~input_layer[1074]),
      .c(~input_layer[1154]),
      .d(input_layer[553]),
      .e(~input_layer[61]),
      .f(~input_layer[163]),
      .y(Y[1008]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_315 for neuron1009_1
  function_315 neuron1009_1 (
      .a(~input_layer[1166]),
      .b(~input_layer[1003]),
      .c(input_layer[566]),
      .d(input_layer[143]),
      .e(input_layer[768]),
      .f(input_layer[397]),
      .y(Y[1009]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1010_1
  function_10 neuron1010_1 (
      .a(~input_layer[799]),
      .b(input_layer[556]),
      .c(input_layer[1150]),
      .d(~input_layer[440]),
      .e(input_layer[527]),
      .f(~input_layer[1230]),
      .y(Y[1010]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_316 for neuron1011_1
  function_316 neuron1011_1 (
      .a(~input_layer[1159]),
      .b(input_layer[1034]),
      .c(~input_layer[1337]),
      .d(~input_layer[925]),
      .e(input_layer[1554]),
      .f(~input_layer[1174]),
      .y(Y[1011]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1012_1
  function_39 neuron1012_1 (
      .a(~input_layer[1137]),
      .b(input_layer[440]),
      .c(~input_layer[358]),
      .y(Y[1012]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1013_1
  function_78 neuron1013_1 (
      .a(~input_layer[425]),
      .b(~input_layer[1078]),
      .c(input_layer[639]),
      .d(input_layer[596]),
      .e(input_layer[673]),
      .f(input_layer[282]),
      .y(Y[1013]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron1014_1
  function_290 neuron1014_1 (
      .a(~input_layer[604]),
      .b(input_layer[1037]),
      .c(~input_layer[1323]),
      .d(~input_layer[778]),
      .e(~input_layer[281]),
      .f(input_layer[1285]),
      .y(Y[1014]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1015_1
  function_5 neuron1015_1 (
      .a(~input_layer[307]),
      .b(~input_layer[1140]),
      .c(~input_layer[265]),
      .d(input_layer[625]),
      .e(~input_layer[433]),
      .f(input_layer[577]),
      .y(Y[1015]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1016_1
  function_0 neuron1016_1 (
      .a(~input_layer[646]),
      .b(~input_layer[1333]),
      .c(input_layer[1197]),
      .d(~input_layer[1378]),
      .e(~input_layer[1124]),
      .y(Y[1016]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1017_1
  function_0 neuron1017_1 (
      .a(~input_layer[187]),
      .b(~input_layer[409]),
      .c(~input_layer[958]),
      .d(input_layer[91]),
      .e(~input_layer[601]),
      .y(Y[1017]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1018_1
  function_19 neuron1018_1 (
      .a(input_layer[465]),
      .b(~input_layer[773]),
      .c(~input_layer[1282]),
      .d(~input_layer[286]),
      .y(Y[1018]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron1019_1
  function_70 neuron1019_1 (
      .a(~input_layer[736]),
      .b(~input_layer[400]),
      .c(input_layer[1050]),
      .d(input_layer[86]),
      .e(~input_layer[295]),
      .f(~input_layer[44]),
      .y(Y[1019]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_317 for neuron1020_1
  function_317 neuron1020_1 (
      .a(~input_layer[1187]),
      .b(input_layer[1433]),
      .c(input_layer[215]),
      .d(input_layer[612]),
      .e(~input_layer[705]),
      .f(input_layer[145]),
      .y(Y[1020]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1021] = 1'b0;

  // instantiate function_265 for neuron1022_1
  function_265 neuron1022_1 (
      .a(input_layer[495]),
      .b(~input_layer[867]),
      .c(~input_layer[546]),
      .d(input_layer[691]),
      .e(~input_layer[122]),
      .f(input_layer[477]),
      .y(Y[1022]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1023_1
  function_24 neuron1023_1 (
      .a(~input_layer[440]),
      .b(input_layer[703]),
      .c(~input_layer[652]),
      .y(Y[1023]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron1024_1
  function_145 neuron1024_1 (
      .a(input_layer[320]),
      .b(~input_layer[420]),
      .c(~input_layer[513]),
      .d(input_layer[1153]),
      .e(~input_layer[416]),
      .y(Y[1024]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1025_1
  function_29 neuron1025_1 (
      .a(~input_layer[430]),
      .b(input_layer[205]),
      .y(Y[1025]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_318 for neuron1026_1
  function_318 neuron1026_1 (
      .a(input_layer[1370]),
      .b(input_layer[1204]),
      .c(~input_layer[771]),
      .d(~input_layer[147]),
      .e(~input_layer[734]),
      .f(input_layer[1211]),
      .y(Y[1026]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1027_1
  function_135 neuron1027_1 (
      .a(input_layer[1484]),
      .b(input_layer[1480]),
      .c(~input_layer[136]),
      .d(input_layer[637]),
      .e(input_layer[1502]),
      .y(Y[1027]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1028_1
  function_8 neuron1028_1 (
      .a(input_layer[522]),
      .b(input_layer[1226]),
      .c(~input_layer[343]),
      .d(input_layer[158]),
      .y(Y[1028]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_2 for neuron1029_1
  function_2 neuron1029_1 (
      .a(input_layer[946]),
      .b(input_layer[478]),
      .c(~input_layer[689]),
      .d(~input_layer[1309]),
      .e(input_layer[723]),
      .f(~input_layer[1258]),
      .y(Y[1029]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1030_1
  function_113 neuron1030_1 (
      .a(input_layer[701]),
      .b(~input_layer[1537]),
      .c(input_layer[948]),
      .d(~input_layer[543]),
      .e(input_layer[1496]),
      .y(Y[1030]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1031_1
  function_55 neuron1031_1 (
      .a(~input_layer[693]),
      .b(~input_layer[718]),
      .c(~input_layer[820]),
      .d(~input_layer[131]),
      .e(~input_layer[685]),
      .y(Y[1031]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_278 for neuron1032_1
  function_278 neuron1032_1 (
      .a(input_layer[998]),
      .b(~input_layer[624]),
      .c(input_layer[238]),
      .d(input_layer[293]),
      .e(~input_layer[508]),
      .y(Y[1032]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1033_1
  function_28 neuron1033_1 (
      .a(~input_layer[401]),
      .b(~input_layer[371]),
      .c(~input_layer[620]),
      .d(~input_layer[1060]),
      .e(~input_layer[1447]),
      .f(~input_layer[1229]),
      .y(Y[1033]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1034_1
  function_27 neuron1034_1 (
      .a(~input_layer[1106]),
      .b(~input_layer[370]),
      .c(~input_layer[204]),
      .y(Y[1034]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1035_1
  function_42 neuron1035_1 (
      .a(input_layer[188]),
      .b(input_layer[240]),
      .c(input_layer[272]),
      .d(input_layer[177]),
      .y(Y[1035]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron1036_1
  function_96 neuron1036_1 (
      .a(input_layer[1381]),
      .b(input_layer[1264]),
      .c(~input_layer[1466]),
      .d(~input_layer[777]),
      .y(Y[1036]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1037_1
  function_319 neuron1037_1 (
      .a(input_layer[909]),
      .b(~input_layer[1208]),
      .c(input_layer[798]),
      .d(~input_layer[585]),
      .e(~input_layer[450]),
      .f(input_layer[436]),
      .y(Y[1037]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_320 for neuron1038_1
  function_320 neuron1038_1 (
      .a(input_layer[1057]),
      .b(~input_layer[748]),
      .c(~input_layer[131]),
      .d(~input_layer[864]),
      .e(input_layer[879]),
      .f(input_layer[30]),
      .y(Y[1038]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_321 for neuron1039_1
  function_321 neuron1039_1 (
      .a(input_layer[292]),
      .b(~input_layer[637]),
      .c(input_layer[131]),
      .d(input_layer[467]),
      .e(input_layer[308]),
      .f(input_layer[1393]),
      .y(Y[1039]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1040_1
  function_24 neuron1040_1 (
      .a(~input_layer[487]),
      .b(~input_layer[592]),
      .c(input_layer[1082]),
      .y(Y[1040]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1041_1
  function_42 neuron1041_1 (
      .a(input_layer[191]),
      .b(input_layer[1296]),
      .c(input_layer[1364]),
      .d(input_layer[623]),
      .y(Y[1041]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1042_1
  function_5 neuron1042_1 (
      .a(~input_layer[425]),
      .b(~input_layer[1227]),
      .c(~input_layer[531]),
      .d(~input_layer[340]),
      .e(input_layer[1094]),
      .f(~input_layer[161]),
      .y(Y[1042]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1043] = 1'b0;

  // instantiate function_67 for neuron1044_1
  function_67 neuron1044_1 (
      .a(~input_layer[768]),
      .b(~input_layer[399]),
      .c(~input_layer[1408]),
      .d(~input_layer[650]),
      .e(input_layer[1191]),
      .y(Y[1044]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_322 for neuron1045_1
  function_322 neuron1045_1 (
      .a(input_layer[1017]),
      .b(~input_layer[803]),
      .c(input_layer[833]),
      .d(~input_layer[1414]),
      .e(input_layer[937]),
      .f(input_layer[363]),
      .y(Y[1045]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_323 for neuron1046_1
  function_323 neuron1046_1 (
      .a(~input_layer[1320]),
      .b(input_layer[1081]),
      .c(input_layer[264]),
      .d(input_layer[208]),
      .e(input_layer[367]),
      .f(input_layer[722]),
      .y(Y[1046]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1047_1
  function_37 neuron1047_1 (
      .a(input_layer[685]),
      .b(input_layer[1482]),
      .c(~input_layer[301]),
      .d(~input_layer[1339]),
      .e(input_layer[955]),
      .f(input_layer[160]),
      .y(Y[1047]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1048_1
  function_27 neuron1048_1 (
      .a(~input_layer[417]),
      .b(~input_layer[1297]),
      .c(~input_layer[1236]),
      .y(Y[1048]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1049_1
  function_107 neuron1049_1 (
      .a(~input_layer[754]),
      .b(~input_layer[979]),
      .c(~input_layer[1157]),
      .d(input_layer[456]),
      .e(~input_layer[804]),
      .y(Y[1049]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron1050_1
  function_65 neuron1050_1 (
      .a(input_layer[703]),
      .b(~input_layer[1092]),
      .c(input_layer[289]),
      .d(input_layer[992]),
      .e(~input_layer[334]),
      .f(~input_layer[103]),
      .y(Y[1050]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1051_1
  function_97 neuron1051_1 (
      .a(~input_layer[1165]),
      .b(~input_layer[893]),
      .c(~input_layer[564]),
      .d(input_layer[95]),
      .e(input_layer[667]),
      .y(Y[1051]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1052_1
  function_31 neuron1052_1 (
      .a(input_layer[1136]),
      .b(~input_layer[1547]),
      .c(~input_layer[512]),
      .d(input_layer[1440]),
      .y(Y[1052]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1053_1
  function_42 neuron1053_1 (
      .a(input_layer[995]),
      .b(input_layer[1047]),
      .c(input_layer[357]),
      .d(input_layer[1181]),
      .y(Y[1053]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_324 for neuron1054_1
  function_324 neuron1054_1 (
      .a(~input_layer[883]),
      .b(input_layer[576]),
      .c(~input_layer[1074]),
      .d(input_layer[1393]),
      .e(input_layer[1406]),
      .y(Y[1054]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1055_1
  function_29 neuron1055_1 (
      .a(~input_layer[246]),
      .b(input_layer[522]),
      .y(Y[1055]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1056_1
  function_0 neuron1056_1 (
      .a(~input_layer[831]),
      .b(~input_layer[916]),
      .c(~input_layer[779]),
      .d(input_layer[366]),
      .e(~input_layer[1009]),
      .y(Y[1056]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1057_1
  function_24 neuron1057_1 (
      .a(~input_layer[878]),
      .b(input_layer[1315]),
      .c(input_layer[1314]),
      .y(Y[1057]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1058_1
  function_19 neuron1058_1 (
      .a(~input_layer[259]),
      .b(~input_layer[212]),
      .c(~input_layer[93]),
      .d(input_layer[618]),
      .y(Y[1058]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_291 for neuron1059_1
  function_291 neuron1059_1 (
      .a(input_layer[263]),
      .b(input_layer[996]),
      .c(~input_layer[1388]),
      .d(input_layer[588]),
      .e(~input_layer[861]),
      .y(Y[1059]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_305 for neuron1060_1
  function_305 neuron1060_1 (
      .a(~input_layer[297]),
      .b(input_layer[542]),
      .c(input_layer[677]),
      .d(~input_layer[1351]),
      .e(~input_layer[285]),
      .y(Y[1060]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1061_1
  function_181 neuron1061_1 (
      .a(input_layer[1029]),
      .b(~input_layer[454]),
      .c(input_layer[1324]),
      .d(input_layer[199]),
      .e(~input_layer[1365]),
      .y(Y[1061]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1062_1
  function_42 neuron1062_1 (
      .a(input_layer[779]),
      .b(input_layer[645]),
      .c(input_layer[1254]),
      .d(input_layer[450]),
      .y(Y[1062]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1063_1
  function_29 neuron1063_1 (
      .a(~input_layer[150]),
      .b(input_layer[868]),
      .y(Y[1063]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1064_1
  function_29 neuron1064_1 (
      .a(input_layer[698]),
      .b(~input_layer[625]),
      .y(Y[1064]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_325 for neuron1065_1
  function_325 neuron1065_1 (
      .a(~input_layer[1440]),
      .b(~input_layer[710]),
      .c(input_layer[1161]),
      .d(input_layer[179]),
      .e(~input_layer[712]),
      .f(input_layer[1273]),
      .y(Y[1065]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_326 for neuron1066_1
  function_326 neuron1066_1 (
      .a(~input_layer[1193]),
      .b(input_layer[411]),
      .c(input_layer[507]),
      .d(~input_layer[419]),
      .e(input_layer[160]),
      .f(~input_layer[667]),
      .y(Y[1066]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_327 for neuron1067_1
  function_327 neuron1067_1 (
      .a(input_layer[793]),
      .b(~input_layer[490]),
      .c(~input_layer[556]),
      .d(input_layer[1122]),
      .e(input_layer[69]),
      .f(input_layer[86]),
      .y(Y[1067]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron1068_1
  function_84 neuron1068_1 (
      .a(~input_layer[1077]),
      .b(~input_layer[948]),
      .c(input_layer[1068]),
      .d(~input_layer[81]),
      .e(input_layer[829]),
      .y(Y[1068]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_328 for neuron1069_1
  function_328 neuron1069_1 (
      .a(~input_layer[1170]),
      .b(~input_layer[358]),
      .c(input_layer[805]),
      .d(input_layer[621]),
      .e(input_layer[94]),
      .f(input_layer[728]),
      .y(Y[1069]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_329 for neuron1070_1
  function_329 neuron1070_1 (
      .a(~input_layer[591]),
      .b(input_layer[684]),
      .c(~input_layer[356]),
      .d(input_layer[850]),
      .e(input_layer[1229]),
      .f(~input_layer[38]),
      .y(Y[1070]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_245 for neuron1071_1
  function_245 neuron1071_1 (
      .a(~input_layer[349]),
      .b(input_layer[1485]),
      .c(input_layer[583]),
      .d(input_layer[97]),
      .e(~input_layer[598]),
      .f(input_layer[779]),
      .y(Y[1071]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1072_1
  function_123 neuron1072_1 (
      .a(input_layer[1372]),
      .b(~input_layer[915]),
      .c(~input_layer[242]),
      .d(~input_layer[564]),
      .y(Y[1072]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1073_1
  function_330 neuron1073_1 (
      .a(~input_layer[690]),
      .b(~input_layer[331]),
      .c(input_layer[398]),
      .d(input_layer[1217]),
      .e(input_layer[1393]),
      .y(Y[1073]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_269 for neuron1074_1
  function_269 neuron1074_1 (
      .a(input_layer[483]),
      .b(input_layer[1014]),
      .c(input_layer[327]),
      .d(input_layer[1012]),
      .e(~input_layer[1093]),
      .f(~input_layer[217]),
      .y(Y[1074]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1075_1
  function_16 neuron1075_1 (
      .a(input_layer[131]),
      .b(~input_layer[657]),
      .y(Y[1075]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1076_1
  function_149 neuron1076_1 (
      .a(input_layer[1258]),
      .b(~input_layer[1333]),
      .c(input_layer[628]),
      .d(~input_layer[882]),
      .y(Y[1076]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1077_1
  function_16 neuron1077_1 (
      .a(~input_layer[813]),
      .b(input_layer[211]),
      .y(Y[1077]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1078_1
  function_76 neuron1078_1 (
      .a(input_layer[1057]),
      .b(input_layer[554]),
      .c(input_layer[79]),
      .d(input_layer[1535]),
      .e(~input_layer[416]),
      .f(~input_layer[414]),
      .y(Y[1078]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1079_1
  function_106 neuron1079_1 (
      .a(input_layer[1165]),
      .b(input_layer[127]),
      .c(input_layer[1252]),
      .d(~input_layer[978]),
      .y(Y[1079]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1080_1
  function_35 neuron1080_1 (
      .a(~input_layer[405]),
      .b(~input_layer[1212]),
      .c(input_layer[485]),
      .d(~input_layer[502]),
      .e(~input_layer[100]),
      .y(Y[1080]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1081_1
  function_95 neuron1081_1 (
      .a(~input_layer[1189]),
      .b(input_layer[1429]),
      .c(input_layer[476]),
      .d(input_layer[182]),
      .y(Y[1081]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1082_1
  function_26 neuron1082_1 (
      .a(input_layer[1335]),
      .y(Y[1082]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_331 for neuron1083_1
  function_331 neuron1083_1 (
      .a(input_layer[459]),
      .b(~input_layer[81]),
      .c(input_layer[1530]),
      .d(~input_layer[219]),
      .e(input_layer[1524]),
      .f(~input_layer[816]),
      .y(Y[1083]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1084_1
  function_148 neuron1084_1 (
      .a(input_layer[421]),
      .b(input_layer[1302]),
      .c(~input_layer[651]),
      .d(input_layer[101]),
      .e(~input_layer[969]),
      .f(input_layer[43]),
      .y(Y[1084]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1085_1
  function_5 neuron1085_1 (
      .a(~input_layer[417]),
      .b(~input_layer[304]),
      .c(~input_layer[1309]),
      .d(input_layer[866]),
      .e(input_layer[939]),
      .f(~input_layer[995]),
      .y(Y[1085]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1086_1
  function_17 neuron1086_1 (
      .a(input_layer[417]),
      .b(~input_layer[585]),
      .c(input_layer[185]),
      .y(Y[1086]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron1087_1
  function_155 neuron1087_1 (
      .a(~input_layer[1157]),
      .b(~input_layer[1330]),
      .c(~input_layer[389]),
      .d(~input_layer[910]),
      .e(input_layer[156]),
      .f(~input_layer[1405]),
      .y(Y[1087]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1088_1
  function_17 neuron1088_1 (
      .a(input_layer[407]),
      .b(input_layer[581]),
      .c(input_layer[322]),
      .y(Y[1088]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1089_1
  function_126 neuron1089_1 (
      .a(~input_layer[1081]),
      .b(~input_layer[1103]),
      .c(input_layer[512]),
      .d(~input_layer[153]),
      .e(~input_layer[241]),
      .y(Y[1089]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1090_1
  function_0 neuron1090_1 (
      .a(~input_layer[1472]),
      .b(~input_layer[130]),
      .c(~input_layer[182]),
      .d(~input_layer[535]),
      .e(input_layer[1188]),
      .y(Y[1090]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1091_1
  function_16 neuron1091_1 (
      .a(input_layer[1003]),
      .b(input_layer[1192]),
      .y(Y[1091]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1092_1
  function_120 neuron1092_1 (
      .a(input_layer[929]),
      .b(input_layer[200]),
      .c(~input_layer[964]),
      .d(input_layer[1394]),
      .e(~input_layer[274]),
      .y(Y[1092]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1093_1
  function_172 neuron1093_1 (
      .a(~input_layer[312]),
      .b(~input_layer[499]),
      .c(~input_layer[1130]),
      .d(~input_layer[436]),
      .e(~input_layer[1295]),
      .f(input_layer[797]),
      .y(Y[1093]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1094_1
  function_135 neuron1094_1 (
      .a(~input_layer[966]),
      .b(input_layer[1161]),
      .c(input_layer[949]),
      .d(input_layer[390]),
      .e(input_layer[1178]),
      .y(Y[1094]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1095_1
  function_271 neuron1095_1 (
      .a(~input_layer[1431]),
      .b(input_layer[1015]),
      .c(input_layer[127]),
      .d(input_layer[1319]),
      .e(input_layer[1311]),
      .y(Y[1095]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1096_1
  function_126 neuron1096_1 (
      .a(~input_layer[523]),
      .b(input_layer[252]),
      .c(~input_layer[823]),
      .d(input_layer[869]),
      .e(~input_layer[265]),
      .y(Y[1096]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1097_1
  function_54 neuron1097_1 (
      .a(input_layer[191]),
      .b(~input_layer[600]),
      .c(input_layer[212]),
      .d(~input_layer[904]),
      .e(input_layer[1556]),
      .f(input_layer[361]),
      .y(Y[1097]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_332 for neuron1098_1
  function_332 neuron1098_1 (
      .a(~input_layer[1154]),
      .b(input_layer[1537]),
      .c(~input_layer[689]),
      .d(input_layer[424]),
      .e(~input_layer[151]),
      .f(~input_layer[557]),
      .y(Y[1098]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1099_1
  function_162 neuron1099_1 (
      .a(input_layer[1001]),
      .b(input_layer[1162]),
      .c(~input_layer[325]),
      .d(input_layer[1134]),
      .e(~input_layer[1390]),
      .f(~input_layer[479]),
      .y(Y[1099]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1100_1
  function_298 neuron1100_1 (
      .a(~input_layer[1494]),
      .b(~input_layer[425]),
      .c(~input_layer[333]),
      .d(~input_layer[817]),
      .e(input_layer[969]),
      .f(~input_layer[1211]),
      .y(Y[1100]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1101_1
  function_5 neuron1101_1 (
      .a(~input_layer[1278]),
      .b(~input_layer[859]),
      .c(~input_layer[189]),
      .d(input_layer[379]),
      .e(input_layer[1093]),
      .f(input_layer[232]),
      .y(Y[1101]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1102_1
  function_106 neuron1102_1 (
      .a(input_layer[915]),
      .b(input_layer[886]),
      .c(input_layer[485]),
      .d(input_layer[937]),
      .y(Y[1102]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1103_1
  function_39 neuron1103_1 (
      .a(~input_layer[855]),
      .b(input_layer[1380]),
      .c(~input_layer[914]),
      .y(Y[1103]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1104_1
  function_46 neuron1104_1 (
      .a(input_layer[1070]),
      .b(~input_layer[1260]),
      .c(input_layer[1125]),
      .d(input_layer[1167]),
      .e(~input_layer[622]),
      .y(Y[1104]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1105_1
  function_128 neuron1105_1 (
      .a(~input_layer[1440]),
      .b(input_layer[1160]),
      .c(input_layer[568]),
      .d(~input_layer[1376]),
      .y(Y[1105]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_333 for neuron1106_1
  function_333 neuron1106_1 (
      .a(~input_layer[1184]),
      .b(input_layer[153]),
      .c(input_layer[156]),
      .d(input_layer[1027]),
      .e(~input_layer[869]),
      .f(~input_layer[479]),
      .y(Y[1106]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1107_1
  function_76 neuron1107_1 (
      .a(input_layer[612]),
      .b(input_layer[326]),
      .c(input_layer[725]),
      .d(input_layer[562]),
      .e(~input_layer[473]),
      .f(input_layer[24]),
      .y(Y[1107]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1108_1
  function_8 neuron1108_1 (
      .a(input_layer[978]),
      .b(input_layer[454]),
      .c(~input_layer[372]),
      .d(input_layer[96]),
      .y(Y[1108]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1109_1
  function_27 neuron1109_1 (
      .a(~input_layer[1480]),
      .b(~input_layer[753]),
      .c(~input_layer[886]),
      .y(Y[1109]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1110_1
  function_24 neuron1110_1 (
      .a(~input_layer[1095]),
      .b(~input_layer[158]),
      .c(input_layer[1473]),
      .y(Y[1110]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron1111_1
  function_121 neuron1111_1 (
      .a(input_layer[1319]),
      .b(input_layer[346]),
      .c(input_layer[1530]),
      .d(~input_layer[1052]),
      .e(~input_layer[853]),
      .y(Y[1111]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron1112_1
  function_69 neuron1112_1 (
      .a(input_layer[645]),
      .b(~input_layer[1089]),
      .c(~input_layer[941]),
      .d(~input_layer[1122]),
      .e(input_layer[1523]),
      .f(input_layer[1342]),
      .y(Y[1112]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1113_1
  function_334 neuron1113_1 (
      .a(~input_layer[661]),
      .b(input_layer[1049]),
      .c(input_layer[1158]),
      .d(input_layer[1139]),
      .e(~input_layer[1368]),
      .y(Y[1113]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_335 for neuron1114_1
  function_335 neuron1114_1 (
      .a(~input_layer[1483]),
      .b(~input_layer[877]),
      .c(~input_layer[623]),
      .d(input_layer[1263]),
      .e(input_layer[447]),
      .f(input_layer[934]),
      .y(Y[1114]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1115_1
  function_126 neuron1115_1 (
      .a(~input_layer[1161]),
      .b(~input_layer[610]),
      .c(~input_layer[1280]),
      .d(~input_layer[751]),
      .e(input_layer[823]),
      .y(Y[1115]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1116_1
  function_25 neuron1116_1 (
      .a(~input_layer[798]),
      .b(input_layer[514]),
      .c(input_layer[247]),
      .d(input_layer[643]),
      .e(input_layer[609]),
      .y(Y[1116]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron1117_1
  function_36 neuron1117_1 (
      .a(input_layer[1476]),
      .b(input_layer[633]),
      .c(~input_layer[642]),
      .d(input_layer[557]),
      .e(input_layer[1493]),
      .f(input_layer[276]),
      .y(Y[1117]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1118_1
  function_46 neuron1118_1 (
      .a(input_layer[1185]),
      .b(~input_layer[528]),
      .c(input_layer[181]),
      .d(input_layer[1201]),
      .e(input_layer[319]),
      .y(Y[1118]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1119_1
  function_271 neuron1119_1 (
      .a(~input_layer[856]),
      .b(input_layer[701]),
      .c(input_layer[567]),
      .d(input_layer[1001]),
      .e(input_layer[27]),
      .y(Y[1119]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1120_1
  function_27 neuron1120_1 (
      .a(~input_layer[212]),
      .b(~input_layer[1239]),
      .c(input_layer[1256]),
      .y(Y[1120]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1121_1
  function_17 neuron1121_1 (
      .a(input_layer[456]),
      .b(~input_layer[1314]),
      .c(~input_layer[1154]),
      .y(Y[1121]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_15 for neuron1122_1
  function_15 neuron1122_1 (
      .a(input_layer[834]),
      .b(input_layer[207]),
      .c(~input_layer[930]),
      .d(input_layer[1527]),
      .e(input_layer[518]),
      .f(~input_layer[1011]),
      .y(Y[1122]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1123_1
  function_19 neuron1123_1 (
      .a(~input_layer[207]),
      .b(~input_layer[1210]),
      .c(~input_layer[83]),
      .d(input_layer[1531]),
      .y(Y[1123]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_336 for neuron1124_1
  function_336 neuron1124_1 (
      .a(~input_layer[1377]),
      .b(input_layer[1164]),
      .c(~input_layer[645]),
      .d(input_layer[316]),
      .e(~input_layer[1449]),
      .f(~input_layer[396]),
      .y(Y[1124]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1125_1
  function_95 neuron1125_1 (
      .a(~input_layer[907]),
      .b(input_layer[1540]),
      .c(input_layer[668]),
      .d(input_layer[27]),
      .y(Y[1125]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1126_1
  function_11 neuron1126_1 (
      .a(~input_layer[441]),
      .b(input_layer[871]),
      .c(~input_layer[689]),
      .d(input_layer[864]),
      .y(Y[1126]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1127] = 1'b1;

  // instantiate function_19 for neuron1128_1
  function_19 neuron1128_1 (
      .a(~input_layer[199]),
      .b(input_layer[922]),
      .c(~input_layer[929]),
      .d(~input_layer[1389]),
      .y(Y[1128]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1129_1
  function_30 neuron1129_1 (
      .a(input_layer[1372]),
      .b(~input_layer[931]),
      .c(input_layer[151]),
      .d(input_layer[826]),
      .y(Y[1129]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1130_1
  function_26 neuron1130_1 (
      .a(input_layer[700]),
      .y(Y[1130]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_337 for neuron1131_1
  function_337 neuron1131_1 (
      .a(~input_layer[741]),
      .b(input_layer[1115]),
      .c(~input_layer[1440]),
      .d(input_layer[1158]),
      .e(input_layer[461]),
      .f(~input_layer[1500]),
      .y(Y[1131]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1132_1
  function_95 neuron1132_1 (
      .a(~input_layer[194]),
      .b(input_layer[387]),
      .c(input_layer[631]),
      .d(input_layer[684]),
      .y(Y[1132]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1133_1
  function_39 neuron1133_1 (
      .a(~input_layer[1217]),
      .b(input_layer[1491]),
      .c(~input_layer[1045]),
      .y(Y[1133]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_338 for neuron1134_1
  function_338 neuron1134_1 (
      .a(input_layer[428]),
      .b(input_layer[484]),
      .c(input_layer[1191]),
      .d(~input_layer[1351]),
      .e(~input_layer[876]),
      .f(input_layer[1163]),
      .y(Y[1134]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1135_1
  function_45 neuron1135_1 (
      .a(input_layer[1540]),
      .b(input_layer[407]),
      .c(input_layer[453]),
      .d(~input_layer[856]),
      .e(input_layer[1528]),
      .f(input_layer[267]),
      .y(Y[1135]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_339 for neuron1136_1
  function_339 neuron1136_1 (
      .a(~input_layer[692]),
      .b(input_layer[813]),
      .c(~input_layer[1266]),
      .d(input_layer[530]),
      .e(input_layer[1147]),
      .f(input_layer[985]),
      .y(Y[1136]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1137_1
  function_3 neuron1137_1 (
      .a(~input_layer[369]),
      .b(~input_layer[1076]),
      .c(~input_layer[259]),
      .d(~input_layer[348]),
      .y(Y[1137]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1138_1
  function_123 neuron1138_1 (
      .a(input_layer[1142]),
      .b(~input_layer[149]),
      .c(input_layer[626]),
      .d(input_layer[1470]),
      .y(Y[1138]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_340 for neuron1139_1
  function_340 neuron1139_1 (
      .a(~input_layer[1242]),
      .b(~input_layer[1265]),
      .c(input_layer[603]),
      .d(input_layer[96]),
      .e(input_layer[177]),
      .f(~input_layer[780]),
      .y(Y[1139]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1140_1
  function_3 neuron1140_1 (
      .a(~input_layer[1105]),
      .b(~input_layer[738]),
      .c(~input_layer[1532]),
      .d(input_layer[321]),
      .y(Y[1140]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1141_1
  function_214 neuron1141_1 (
      .a(input_layer[1485]),
      .b(~input_layer[378]),
      .c(input_layer[1013]),
      .d(input_layer[845]),
      .e(input_layer[136]),
      .f(input_layer[123]),
      .y(Y[1141]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1142_1
  function_55 neuron1142_1 (
      .a(~input_layer[807]),
      .b(~input_layer[148]),
      .c(~input_layer[691]),
      .d(~input_layer[851]),
      .e(input_layer[1319]),
      .y(Y[1142]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1143_1
  function_67 neuron1143_1 (
      .a(~input_layer[1485]),
      .b(~input_layer[1195]),
      .c(~input_layer[1352]),
      .d(~input_layer[1547]),
      .e(~input_layer[429]),
      .y(Y[1143]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1144_1
  function_27 neuron1144_1 (
      .a(~input_layer[481]),
      .b(~input_layer[405]),
      .c(~input_layer[205]),
      .y(Y[1144]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1145_1
  function_55 neuron1145_1 (
      .a(~input_layer[381]),
      .b(~input_layer[778]),
      .c(~input_layer[1393]),
      .d(input_layer[125]),
      .e(input_layer[79]),
      .y(Y[1145]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1146_1
  function_100 neuron1146_1 (
      .a(~input_layer[136]),
      .b(~input_layer[1171]),
      .c(~input_layer[858]),
      .d(input_layer[1431]),
      .e(~input_layer[95]),
      .f(input_layer[786]),
      .y(Y[1146]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1147_1
  function_55 neuron1147_1 (
      .a(~input_layer[243]),
      .b(~input_layer[466]),
      .c(~input_layer[414]),
      .d(~input_layer[720]),
      .e(input_layer[156]),
      .y(Y[1147]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1148_1
  function_27 neuron1148_1 (
      .a(~input_layer[301]),
      .b(~input_layer[923]),
      .c(~input_layer[293]),
      .y(Y[1148]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_341 for neuron1149_1
  function_341 neuron1149_1 (
      .a(~input_layer[1086]),
      .b(input_layer[1417]),
      .c(input_layer[1415]),
      .d(~input_layer[999]),
      .e(~input_layer[1252]),
      .f(~input_layer[918]),
      .y(Y[1149]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1150_1
  function_126 neuron1150_1 (
      .a(input_layer[652]),
      .b(~input_layer[1085]),
      .c(~input_layer[1392]),
      .d(~input_layer[1154]),
      .e(~input_layer[1257]),
      .y(Y[1150]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1151_1
  function_42 neuron1151_1 (
      .a(input_layer[1171]),
      .b(input_layer[201]),
      .c(input_layer[1486]),
      .d(input_layer[1229]),
      .y(Y[1151]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1152_1
  function_17 neuron1152_1 (
      .a(input_layer[1143]),
      .b(input_layer[1226]),
      .c(input_layer[126]),
      .y(Y[1152]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1153_1
  function_26 neuron1153_1 (
      .a(~input_layer[983]),
      .y(Y[1153]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1154_1
  function_16 neuron1154_1 (
      .a(input_layer[534]),
      .b(~input_layer[798]),
      .y(Y[1154]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1155_1
  function_78 neuron1155_1 (
      .a(~input_layer[143]),
      .b(~input_layer[591]),
      .c(~input_layer[1001]),
      .d(~input_layer[301]),
      .e(~input_layer[1433]),
      .f(~input_layer[992]),
      .y(Y[1155]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1156_1
  function_0 neuron1156_1 (
      .a(input_layer[441]),
      .b(~input_layer[767]),
      .c(~input_layer[778]),
      .d(~input_layer[623]),
      .e(~input_layer[92]),
      .y(Y[1156]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1157_1
  function_29 neuron1157_1 (
      .a(~input_layer[578]),
      .b(~input_layer[923]),
      .y(Y[1157]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1158_1
  function_29 neuron1158_1 (
      .a(~input_layer[907]),
      .b(input_layer[1262]),
      .y(Y[1158]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_342 for neuron1159_1
  function_342 neuron1159_1 (
      .a(~input_layer[1186]),
      .b(~input_layer[1301]),
      .c(~input_layer[932]),
      .d(input_layer[276]),
      .e(~input_layer[364]),
      .y(Y[1159]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1160_1
  function_26 neuron1160_1 (
      .a(input_layer[796]),
      .y(Y[1160]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_83 for neuron1161_1
  function_83 neuron1161_1 (
      .a(~input_layer[646]),
      .b(input_layer[833]),
      .c(input_layer[885]),
      .d(~input_layer[547]),
      .e(~input_layer[1270]),
      .y(Y[1161]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1162_1
  function_146 neuron1162_1 (
      .a(input_layer[678]),
      .b(input_layer[891]),
      .c(~input_layer[1213]),
      .d(input_layer[618]),
      .e(input_layer[646]),
      .f(input_layer[1066]),
      .y(Y[1162]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1163_1
  function_123 neuron1163_1 (
      .a(input_layer[1430]),
      .b(~input_layer[639]),
      .c(~input_layer[1134]),
      .d(~input_layer[1021]),
      .y(Y[1163]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1164_1
  function_12 neuron1164_1 (
      .a(input_layer[593]),
      .b(~input_layer[322]),
      .c(input_layer[845]),
      .y(Y[1164]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1165_1
  function_29 neuron1165_1 (
      .a(input_layer[299]),
      .b(~input_layer[773]),
      .y(Y[1165]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1166_1
  function_67 neuron1166_1 (
      .a(~input_layer[253]),
      .b(~input_layer[151]),
      .c(~input_layer[366]),
      .d(~input_layer[1159]),
      .e(~input_layer[1047]),
      .y(Y[1166]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_343 for neuron1167_1
  function_343 neuron1167_1 (
      .a(input_layer[330]),
      .b(~input_layer[1496]),
      .c(~input_layer[480]),
      .d(input_layer[638]),
      .e(~input_layer[1117]),
      .f(~input_layer[1123]),
      .y(Y[1167]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1168_1
  function_42 neuron1168_1 (
      .a(input_layer[184]),
      .b(~input_layer[1028]),
      .c(input_layer[183]),
      .d(input_layer[1068]),
      .y(Y[1168]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1169_1
  function_214 neuron1169_1 (
      .a(input_layer[133]),
      .b(input_layer[1301]),
      .c(input_layer[990]),
      .d(input_layer[74]),
      .e(~input_layer[883]),
      .f(input_layer[2]),
      .y(Y[1169]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1170_1
  function_78 neuron1170_1 (
      .a(~input_layer[1279]),
      .b(~input_layer[330]),
      .c(input_layer[515]),
      .d(~input_layer[776]),
      .e(~input_layer[1337]),
      .f(~input_layer[65]),
      .y(Y[1170]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1171_1
  function_27 neuron1171_1 (
      .a(input_layer[422]),
      .b(~input_layer[998]),
      .c(~input_layer[1351]),
      .y(Y[1171]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1172] = 1'b0;

  // instantiate function_128 for neuron1173_1
  function_128 neuron1173_1 (
      .a(~input_layer[799]),
      .b(input_layer[1105]),
      .c(input_layer[391]),
      .d(input_layer[255]),
      .y(Y[1173]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1174_1
  function_8 neuron1174_1 (
      .a(input_layer[694]),
      .b(input_layer[518]),
      .c(input_layer[797]),
      .d(input_layer[1227]),
      .y(Y[1174]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1175_1
  function_27 neuron1175_1 (
      .a(~input_layer[1159]),
      .b(~input_layer[1103]),
      .c(input_layer[462]),
      .y(Y[1175]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1176_1
  function_100 neuron1176_1 (
      .a(~input_layer[1315]),
      .b(~input_layer[739]),
      .c(~input_layer[681]),
      .d(input_layer[862]),
      .e(~input_layer[456]),
      .f(input_layer[319]),
      .y(Y[1176]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_237 for neuron1177_1
  function_237 neuron1177_1 (
      .a(~input_layer[799]),
      .b(input_layer[403]),
      .c(input_layer[949]),
      .d(~input_layer[849]),
      .e(~input_layer[527]),
      .y(Y[1177]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1178_1
  function_97 neuron1178_1 (
      .a(~input_layer[134]),
      .b(~input_layer[313]),
      .c(input_layer[626]),
      .d(~input_layer[1322]),
      .e(~input_layer[94]),
      .y(Y[1178]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1179_1
  function_47 neuron1179_1 (
      .a(input_layer[207]),
      .b(input_layer[1038]),
      .c(input_layer[277]),
      .d(input_layer[262]),
      .e(input_layer[1057]),
      .y(Y[1179]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_304 for neuron1180_1
  function_304 neuron1180_1 (
      .a(~input_layer[200]),
      .b(input_layer[919]),
      .c(input_layer[980]),
      .d(~input_layer[347]),
      .e(~input_layer[1092]),
      .f(~input_layer[840]),
      .y(Y[1180]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1181_1
  function_27 neuron1181_1 (
      .a(~input_layer[202]),
      .b(~input_layer[286]),
      .c(~input_layer[1155]),
      .y(Y[1181]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1182_1
  function_60 neuron1182_1 (
      .a(input_layer[1058]),
      .b(input_layer[240]),
      .c(input_layer[1190]),
      .d(~input_layer[438]),
      .e(input_layer[1100]),
      .y(Y[1182]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1183_1
  function_149 neuron1183_1 (
      .a(~input_layer[646]),
      .b(~input_layer[664]),
      .c(input_layer[1094]),
      .d(~input_layer[704]),
      .y(Y[1183]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1184_1
  function_4 neuron1184_1 (
      .a(~input_layer[656]),
      .b(~input_layer[537]),
      .c(~input_layer[1026]),
      .d(~input_layer[1178]),
      .e(~input_layer[1179]),
      .y(Y[1184]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1185_1
  function_29 neuron1185_1 (
      .a(input_layer[422]),
      .b(~input_layer[1084]),
      .y(Y[1185]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_344 for neuron1186_1
  function_344 neuron1186_1 (
      .a(input_layer[1276]),
      .b(~input_layer[1299]),
      .c(input_layer[91]),
      .d(~input_layer[541]),
      .e(~input_layer[1192]),
      .f(input_layer[223]),
      .y(Y[1186]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_343 for neuron1187_1
  function_343 neuron1187_1 (
      .a(~input_layer[479]),
      .b(~input_layer[716]),
      .c(input_layer[649]),
      .d(~input_layer[1542]),
      .e(input_layer[648]),
      .f(input_layer[1269]),
      .y(Y[1187]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_279 for neuron1188_1
  function_279 neuron1188_1 (
      .a(~input_layer[808]),
      .b(input_layer[1490]),
      .c(input_layer[1484]),
      .d(~input_layer[644]),
      .e(~input_layer[956]),
      .y(Y[1188]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1189_1
  function_8 neuron1189_1 (
      .a(input_layer[1375]),
      .b(input_layer[1278]),
      .c(input_layer[458]),
      .d(input_layer[1472]),
      .y(Y[1189]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1190_1
  function_78 neuron1190_1 (
      .a(~input_layer[1115]),
      .b(~input_layer[856]),
      .c(input_layer[546]),
      .d(~input_layer[844]),
      .e(~input_layer[98]),
      .f(~input_layer[729]),
      .y(Y[1190]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1191_1
  function_67 neuron1191_1 (
      .a(~input_layer[744]),
      .b(~input_layer[350]),
      .c(~input_layer[461]),
      .d(~input_layer[1441]),
      .e(~input_layer[383]),
      .y(Y[1191]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron1192_1
  function_290 neuron1192_1 (
      .a(~input_layer[806]),
      .b(~input_layer[974]),
      .c(~input_layer[1249]),
      .d(input_layer[735]),
      .e(input_layer[1009]),
      .f(input_layer[1502]),
      .y(Y[1192]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1193_1
  function_0 neuron1193_1 (
      .a(~input_layer[1048]),
      .b(~input_layer[130]),
      .c(~input_layer[260]),
      .d(input_layer[520]),
      .e(~input_layer[1259]),
      .y(Y[1193]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_345 for neuron1194_1
  function_345 neuron1194_1 (
      .a(input_layer[1222]),
      .b(input_layer[1436]),
      .c(~input_layer[995]),
      .d(~input_layer[699]),
      .e(input_layer[1489]),
      .f(input_layer[359]),
      .y(Y[1194]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1195_1
  function_17 neuron1195_1 (
      .a(input_layer[486]),
      .b(input_layer[1329]),
      .c(input_layer[1171]),
      .y(Y[1195]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_255 for neuron1196_1
  function_255 neuron1196_1 (
      .a(input_layer[652]),
      .b(~input_layer[836]),
      .c(~input_layer[124]),
      .d(~input_layer[1408]),
      .e(input_layer[243]),
      .y(Y[1196]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1197_1
  function_27 neuron1197_1 (
      .a(~input_layer[981]),
      .b(~input_layer[1436]),
      .c(~input_layer[188]),
      .y(Y[1197]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1198_1
  function_19 neuron1198_1 (
      .a(~input_layer[499]),
      .b(~input_layer[1279]),
      .c(input_layer[1193]),
      .d(input_layer[1305]),
      .y(Y[1198]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1199_1
  function_26 neuron1199_1 (
      .a(input_layer[534]),
      .y(Y[1199]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1200_1
  function_17 neuron1200_1 (
      .a(input_layer[1002]),
      .b(~input_layer[977]),
      .c(input_layer[850]),
      .y(Y[1200]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_346 for neuron1201_1
  function_346 neuron1201_1 (
      .a(input_layer[1489]),
      .b(~input_layer[1193]),
      .c(input_layer[929]),
      .d(~input_layer[332]),
      .e(~input_layer[944]),
      .f(input_layer[119]),
      .y(Y[1201]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_347 for neuron1202_1
  function_347 neuron1202_1 (
      .a(input_layer[1075]),
      .b(input_layer[204]),
      .c(~input_layer[1529]),
      .d(~input_layer[549]),
      .e(~input_layer[738]),
      .f(input_layer[926]),
      .y(Y[1202]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1203_1
  function_47 neuron1203_1 (
      .a(input_layer[1305]),
      .b(input_layer[1388]),
      .c(input_layer[458]),
      .d(input_layer[1413]),
      .e(input_layer[535]),
      .y(Y[1203]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1204_1
  function_67 neuron1204_1 (
      .a(~input_layer[1052]),
      .b(~input_layer[1243]),
      .c(~input_layer[824]),
      .d(~input_layer[386]),
      .e(~input_layer[778]),
      .y(Y[1204]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1205_1
  function_89 neuron1205_1 (
      .a(input_layer[931]),
      .b(input_layer[161]),
      .c(input_layer[834]),
      .d(input_layer[1175]),
      .e(~input_layer[383]),
      .y(Y[1205]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1206_1
  function_146 neuron1206_1 (
      .a(input_layer[583]),
      .b(input_layer[1227]),
      .c(~input_layer[644]),
      .d(input_layer[1004]),
      .e(input_layer[1117]),
      .f(input_layer[1421]),
      .y(Y[1206]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_348 for neuron1207_1
  function_348 neuron1207_1 (
      .a(~input_layer[1133]),
      .b(input_layer[714]),
      .c(input_layer[93]),
      .d(~input_layer[743]),
      .e(~input_layer[359]),
      .f(input_layer[120]),
      .y(Y[1207]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_50 for neuron1208_1
  function_50 neuron1208_1 (
      .a(~input_layer[708]),
      .b(input_layer[1109]),
      .c(~input_layer[571]),
      .d(input_layer[446]),
      .e(input_layer[1335]),
      .f(~input_layer[1385]),
      .y(Y[1208]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1209_1
  function_17 neuron1209_1 (
      .a(input_layer[714]),
      .b(input_layer[706]),
      .c(input_layer[664]),
      .y(Y[1209]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1210_1
  function_17 neuron1210_1 (
      .a(input_layer[1132]),
      .b(input_layer[296]),
      .c(input_layer[314]),
      .y(Y[1210]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1211_1
  function_92 neuron1211_1 (
      .a(input_layer[1497]),
      .b(input_layer[360]),
      .c(input_layer[1538]),
      .d(~input_layer[860]),
      .e(input_layer[642]),
      .f(input_layer[288]),
      .y(Y[1211]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1212_1
  function_47 neuron1212_1 (
      .a(input_layer[1247]),
      .b(input_layer[512]),
      .c(input_layer[156]),
      .d(input_layer[89]),
      .e(input_layer[276]),
      .y(Y[1212]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1213_1
  function_39 neuron1213_1 (
      .a(~input_layer[263]),
      .b(input_layer[1427]),
      .c(~input_layer[938]),
      .y(Y[1213]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1214_1
  function_42 neuron1214_1 (
      .a(~input_layer[474]),
      .b(input_layer[609]),
      .c(input_layer[388]),
      .d(input_layer[403]),
      .y(Y[1214]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_349 for neuron1215_1
  function_349 neuron1215_1 (
      .a(input_layer[1353]),
      .b(~input_layer[743]),
      .c(input_layer[347]),
      .d(input_layer[880]),
      .e(input_layer[511]),
      .y(Y[1215]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron1216_1
  function_131 neuron1216_1 (
      .a(input_layer[501]),
      .b(input_layer[489]),
      .c(~input_layer[186]),
      .d(~input_layer[215]),
      .e(~input_layer[1086]),
      .f(~input_layer[507]),
      .y(Y[1216]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_268 for neuron1217_1
  function_268 neuron1217_1 (
      .a(input_layer[873]),
      .b(~input_layer[387]),
      .c(input_layer[874]),
      .d(~input_layer[217]),
      .e(~input_layer[1319]),
      .f(input_layer[653]),
      .y(Y[1217]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1218_1
  function_91 neuron1218_1 (
      .a(input_layer[1478]),
      .b(~input_layer[1218]),
      .c(input_layer[457]),
      .d(input_layer[502]),
      .e(~input_layer[421]),
      .y(Y[1218]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1219_1
  function_78 neuron1219_1 (
      .a(~input_layer[349]),
      .b(~input_layer[1159]),
      .c(~input_layer[78]),
      .d(~input_layer[275]),
      .e(~input_layer[1406]),
      .f(~input_layer[1453]),
      .y(Y[1219]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_300 for neuron1220_1
  function_300 neuron1220_1 (
      .a(input_layer[1204]),
      .b(input_layer[159]),
      .c(~input_layer[417]),
      .d(input_layer[996]),
      .e(~input_layer[758]),
      .y(Y[1220]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_350 for neuron1221_1
  function_350 neuron1221_1 (
      .a(input_layer[443]),
      .b(~input_layer[1430]),
      .c(~input_layer[1447]),
      .d(input_layer[1206]),
      .e(~input_layer[1477]),
      .y(Y[1221]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1222_1
  function_16 neuron1222_1 (
      .a(input_layer[1364]),
      .b(input_layer[1490]),
      .y(Y[1222]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron1223_1
  function_241 neuron1223_1 (
      .a(input_layer[1470]),
      .b(input_layer[388]),
      .c(input_layer[566]),
      .d(input_layer[666]),
      .e(~input_layer[1233]),
      .f(input_layer[107]),
      .y(Y[1223]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1224_1
  function_26 neuron1224_1 (
      .a(input_layer[1321]),
      .y(Y[1224]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1225_1
  function_128 neuron1225_1 (
      .a(input_layer[1314]),
      .b(~input_layer[219]),
      .c(~input_layer[1397]),
      .d(~input_layer[1457]),
      .y(Y[1225]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_351 for neuron1226_1
  function_351 neuron1226_1 (
      .a(~input_layer[1059]),
      .b(input_layer[1373]),
      .c(~input_layer[738]),
      .d(input_layer[621]),
      .e(~input_layer[1201]),
      .f(~input_layer[1340]),
      .y(Y[1226]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1227_1
  function_231 neuron1227_1 (
      .a(~input_layer[1186]),
      .b(input_layer[1056]),
      .c(~input_layer[752]),
      .d(input_layer[658]),
      .e(input_layer[1551]),
      .f(~input_layer[405]),
      .y(Y[1227]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1228_1
  function_42 neuron1228_1 (
      .a(input_layer[885]),
      .b(input_layer[1417]),
      .c(input_layer[1412]),
      .d(~input_layer[413]),
      .y(Y[1228]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1229_1
  function_27 neuron1229_1 (
      .a(~input_layer[1413]),
      .b(~input_layer[1116]),
      .c(~input_layer[533]),
      .y(Y[1229]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_218 for neuron1230_1
  function_218 neuron1230_1 (
      .a(input_layer[715]),
      .b(~input_layer[298]),
      .c(input_layer[78]),
      .d(~input_layer[420]),
      .e(~input_layer[425]),
      .y(Y[1230]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1231_1
  function_29 neuron1231_1 (
      .a(~input_layer[1371]),
      .b(input_layer[759]),
      .y(Y[1231]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1232_1
  function_4 neuron1232_1 (
      .a(~input_layer[1432]),
      .b(~input_layer[571]),
      .c(input_layer[91]),
      .d(~input_layer[1285]),
      .e(input_layer[1348]),
      .y(Y[1232]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1233_1
  function_4 neuron1233_1 (
      .a(input_layer[920]),
      .b(~input_layer[455]),
      .c(input_layer[1323]),
      .d(~input_layer[340]),
      .e(~input_layer[573]),
      .y(Y[1233]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1234_1
  function_12 neuron1234_1 (
      .a(input_layer[865]),
      .b(~input_layer[1074]),
      .c(input_layer[848]),
      .y(Y[1234]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1235_1
  function_148 neuron1235_1 (
      .a(input_layer[1186]),
      .b(~input_layer[652]),
      .c(input_layer[622]),
      .d(~input_layer[850]),
      .e(input_layer[748]),
      .f(~input_layer[865]),
      .y(Y[1235]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1236_1
  function_90 neuron1236_1 (
      .a(~input_layer[544]),
      .b(~input_layer[1186]),
      .c(~input_layer[1180]),
      .d(input_layer[816]),
      .e(input_layer[814]),
      .y(Y[1236]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_352 for neuron1237_1
  function_352 neuron1237_1 (
      .a(~input_layer[1317]),
      .b(input_layer[1100]),
      .c(input_layer[246]),
      .d(~input_layer[531]),
      .e(~input_layer[424]),
      .f(input_layer[1120]),
      .y(Y[1237]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron1238_1
  function_36 neuron1238_1 (
      .a(input_layer[601]),
      .b(input_layer[987]),
      .c(input_layer[1432]),
      .d(input_layer[686]),
      .e(input_layer[198]),
      .f(~input_layer[1325]),
      .y(Y[1238]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1239_1
  function_42 neuron1239_1 (
      .a(input_layer[1098]),
      .b(input_layer[1104]),
      .c(input_layer[287]),
      .d(~input_layer[1414]),
      .y(Y[1239]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1240_1
  function_42 neuron1240_1 (
      .a(input_layer[1055]),
      .b(~input_layer[700]),
      .c(input_layer[680]),
      .d(input_layer[1168]),
      .y(Y[1240]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_304 for neuron1241_1
  function_304 neuron1241_1 (
      .a(~input_layer[713]),
      .b(input_layer[320]),
      .c(~input_layer[178]),
      .d(input_layer[575]),
      .e(~input_layer[449]),
      .f(~input_layer[9]),
      .y(Y[1241]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_134 for neuron1242_1
  function_134 neuron1242_1 (
      .a(input_layer[457]),
      .b(input_layer[1109]),
      .c(input_layer[1091]),
      .d(input_layer[1170]),
      .e(~input_layer[685]),
      .f(~input_layer[648]),
      .y(Y[1242]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1243_1
  function_67 neuron1243_1 (
      .a(~input_layer[295]),
      .b(~input_layer[1368]),
      .c(~input_layer[1468]),
      .d(~input_layer[1038]),
      .e(~input_layer[846]),
      .y(Y[1243]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1244_1
  function_27 neuron1244_1 (
      .a(~input_layer[1431]),
      .b(~input_layer[314]),
      .c(~input_layer[798]),
      .y(Y[1244]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1245_1
  function_16 neuron1245_1 (
      .a(input_layer[1114]),
      .b(~input_layer[1376]),
      .y(Y[1245]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron1246_1
  function_96 neuron1246_1 (
      .a(~input_layer[636]),
      .b(~input_layer[1379]),
      .c(input_layer[400]),
      .d(~input_layer[655]),
      .y(Y[1246]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_333 for neuron1247_1
  function_333 neuron1247_1 (
      .a(input_layer[248]),
      .b(~input_layer[1410]),
      .c(input_layer[1270]),
      .d(~input_layer[1181]),
      .e(input_layer[1476]),
      .f(input_layer[1548]),
      .y(Y[1247]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1248_1
  function_39 neuron1248_1 (
      .a(~input_layer[1216]),
      .b(input_layer[1013]),
      .c(~input_layer[1187]),
      .y(Y[1248]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1249_1
  function_27 neuron1249_1 (
      .a(~input_layer[563]),
      .b(~input_layer[1091]),
      .c(~input_layer[99]),
      .y(Y[1249]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_353 for neuron1250_1
  function_353 neuron1250_1 (
      .a(input_layer[1260]),
      .b(input_layer[497]),
      .c(~input_layer[1336]),
      .d(~input_layer[992]),
      .e(~input_layer[211]),
      .f(~input_layer[710]),
      .y(Y[1250]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1251_1
  function_0 neuron1251_1 (
      .a(~input_layer[136]),
      .b(~input_layer[1445]),
      .c(~input_layer[735]),
      .d(~input_layer[1017]),
      .e(~input_layer[1179]),
      .y(Y[1251]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1252_1
  function_48 neuron1252_1 (
      .a(input_layer[605]),
      .b(input_layer[402]),
      .c(input_layer[1101]),
      .d(input_layer[1172]),
      .e(~input_layer[1089]),
      .y(Y[1252]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_354 for neuron1253_1
  function_354 neuron1253_1 (
      .a(~input_layer[1314]),
      .b(~input_layer[378]),
      .c(input_layer[1105]),
      .d(input_layer[1082]),
      .e(~input_layer[327]),
      .f(input_layer[317]),
      .y(Y[1253]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_2 for neuron1254_1
  function_2 neuron1254_1 (
      .a(input_layer[1481]),
      .b(~input_layer[1273]),
      .c(input_layer[296]),
      .d(input_layer[513]),
      .e(~input_layer[424]),
      .f(input_layer[617]),
      .y(Y[1254]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1255_1
  function_92 neuron1255_1 (
      .a(input_layer[1436]),
      .b(~input_layer[967]),
      .c(input_layer[329]),
      .d(input_layer[384]),
      .e(input_layer[1554]),
      .f(input_layer[1558]),
      .y(Y[1255]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1256_1
  function_56 neuron1256_1 (
      .a(~input_layer[1304]),
      .b(~input_layer[868]),
      .c(input_layer[1501]),
      .d(input_layer[141]),
      .e(input_layer[231]),
      .y(Y[1256]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1257_1
  function_0 neuron1257_1 (
      .a(~input_layer[130]),
      .b(~input_layer[290]),
      .c(input_layer[744]),
      .d(~input_layer[1528]),
      .e(~input_layer[862]),
      .y(Y[1257]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1258] = 1'b0;

  // instantiate function_3 for neuron1259_1
  function_3 neuron1259_1 (
      .a(~input_layer[832]),
      .b(~input_layer[352]),
      .c(~input_layer[720]),
      .d(~input_layer[1236]),
      .y(Y[1259]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_161 for neuron1260_1
  function_161 neuron1260_1 (
      .a(input_layer[744]),
      .b(~input_layer[681]),
      .c(~input_layer[1056]),
      .d(~input_layer[990]),
      .e(~input_layer[341]),
      .f(input_layer[364]),
      .y(Y[1260]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1261_1
  function_47 neuron1261_1 (
      .a(input_layer[826]),
      .b(input_layer[516]),
      .c(input_layer[525]),
      .d(~input_layer[866]),
      .e(input_layer[1227]),
      .y(Y[1261]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1262_1
  function_42 neuron1262_1 (
      .a(input_layer[986]),
      .b(input_layer[719]),
      .c(input_layer[905]),
      .d(input_layer[890]),
      .y(Y[1262]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_355 for neuron1263_1
  function_355 neuron1263_1 (
      .a(~input_layer[658]),
      .b(~input_layer[130]),
      .c(input_layer[1246]),
      .d(input_layer[1373]),
      .e(input_layer[1212]),
      .f(input_layer[1235]),
      .y(Y[1263]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_184 for neuron1264_1
  function_184 neuron1264_1 (
      .a(~input_layer[1157]),
      .b(input_layer[508]),
      .c(~input_layer[638]),
      .d(~input_layer[1135]),
      .e(input_layer[928]),
      .y(Y[1264]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1265_1
  function_17 neuron1265_1 (
      .a(input_layer[598]),
      .b(input_layer[546]),
      .c(input_layer[569]),
      .y(Y[1265]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1266_1
  function_29 neuron1266_1 (
      .a(~input_layer[192]),
      .b(~input_layer[820]),
      .y(Y[1266]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron1267_1
  function_84 neuron1267_1 (
      .a(~input_layer[741]),
      .b(input_layer[1049]),
      .c(~input_layer[1417]),
      .d(input_layer[1472]),
      .e(input_layer[1311]),
      .y(Y[1267]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1268_1
  function_27 neuron1268_1 (
      .a(~input_layer[914]),
      .b(~input_layer[923]),
      .c(~input_layer[944]),
      .y(Y[1268]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1269_1
  function_26 neuron1269_1 (
      .a(input_layer[643]),
      .y(Y[1269]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_347 for neuron1270_1
  function_347 neuron1270_1 (
      .a(input_layer[1471]),
      .b(input_layer[801]),
      .c(~input_layer[363]),
      .d(~input_layer[1366]),
      .e(input_layer[746]),
      .f(input_layer[266]),
      .y(Y[1270]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_356 for neuron1271_1
  function_356 neuron1271_1 (
      .a(~input_layer[1029]),
      .b(input_layer[1161]),
      .c(input_layer[1311]),
      .d(input_layer[425]),
      .e(~input_layer[821]),
      .f(~input_layer[1488]),
      .y(Y[1271]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_357 for neuron1272_1
  function_357 neuron1272_1 (
      .a(~input_layer[1184]),
      .b(input_layer[580]),
      .c(~input_layer[291]),
      .d(input_layer[557]),
      .e(~input_layer[184]),
      .f(~input_layer[1337]),
      .y(Y[1272]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1273_1
  function_24 neuron1273_1 (
      .a(~input_layer[149]),
      .b(~input_layer[762]),
      .c(input_layer[1205]),
      .y(Y[1273]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_358 for neuron1274_1
  function_358 neuron1274_1 (
      .a(~input_layer[437]),
      .b(~input_layer[431]),
      .c(input_layer[1446]),
      .d(input_layer[778]),
      .e(~input_layer[788]),
      .f(~input_layer[618]),
      .y(Y[1274]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1275_1
  function_87 neuron1275_1 (
      .a(input_layer[597]),
      .b(~input_layer[1264]),
      .c(input_layer[340]),
      .d(input_layer[228]),
      .e(input_layer[162]),
      .y(Y[1275]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1276_1
  function_42 neuron1276_1 (
      .a(input_layer[189]),
      .b(input_layer[998]),
      .c(input_layer[358]),
      .d(input_layer[960]),
      .y(Y[1276]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_359 for neuron1277_1
  function_359 neuron1277_1 (
      .a(input_layer[461]),
      .b(~input_layer[668]),
      .c(input_layer[473]),
      .d(~input_layer[494]),
      .e(input_layer[225]),
      .f(~input_layer[21]),
      .y(Y[1277]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1278_1
  function_39 neuron1278_1 (
      .a(~input_layer[1018]),
      .b(input_layer[748]),
      .c(input_layer[1353]),
      .y(Y[1278]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_360 for neuron1279_1
  function_360 neuron1279_1 (
      .a(input_layer[1163]),
      .b(~input_layer[1068]),
      .c(~input_layer[463]),
      .d(input_layer[1142]),
      .e(~input_layer[618]),
      .y(Y[1279]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1280_1
  function_19 neuron1280_1 (
      .a(~input_layer[203]),
      .b(input_layer[464]),
      .c(~input_layer[1000]),
      .d(input_layer[981]),
      .y(Y[1280]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1281_1
  function_47 neuron1281_1 (
      .a(input_layer[442]),
      .b(input_layer[467]),
      .c(input_layer[1277]),
      .d(input_layer[415]),
      .e(input_layer[564]),
      .y(Y[1281]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1282_1
  function_149 neuron1282_1 (
      .a(~input_layer[706]),
      .b(~input_layer[1378]),
      .c(~input_layer[1446]),
      .d(input_layer[921]),
      .y(Y[1282]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1283_1
  function_27 neuron1283_1 (
      .a(~input_layer[1425]),
      .b(~input_layer[387]),
      .c(input_layer[1033]),
      .y(Y[1283]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1284_1
  function_55 neuron1284_1 (
      .a(input_layer[362]),
      .b(~input_layer[344]),
      .c(~input_layer[94]),
      .d(~input_layer[749]),
      .e(~input_layer[450]),
      .y(Y[1284]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1285_1
  function_67 neuron1285_1 (
      .a(~input_layer[199]),
      .b(~input_layer[1108]),
      .c(~input_layer[240]),
      .d(~input_layer[1499]),
      .e(~input_layer[536]),
      .y(Y[1285]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1286_1
  function_60 neuron1286_1 (
      .a(input_layer[962]),
      .b(~input_layer[1033]),
      .c(input_layer[1116]),
      .d(~input_layer[641]),
      .e(input_layer[616]),
      .y(Y[1286]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1287_1
  function_35 neuron1287_1 (
      .a(~input_layer[1213]),
      .b(~input_layer[1135]),
      .c(~input_layer[1078]),
      .d(~input_layer[700]),
      .e(input_layer[288]),
      .y(Y[1287]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1288_1
  function_172 neuron1288_1 (
      .a(~input_layer[1436]),
      .b(~input_layer[588]),
      .c(~input_layer[1238]),
      .d(~input_layer[1551]),
      .e(~input_layer[559]),
      .f(~input_layer[231]),
      .y(Y[1288]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_361 for neuron1289_1
  function_361 neuron1289_1 (
      .a(~input_layer[1027]),
      .b(input_layer[299]),
      .c(input_layer[620]),
      .d(~input_layer[751]),
      .e(~input_layer[195]),
      .f(~input_layer[1268]),
      .y(Y[1289]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1290_1
  function_20 neuron1290_1 (
      .a(~input_layer[488]),
      .b(~input_layer[1315]),
      .c(input_layer[697]),
      .d(~input_layer[788]),
      .e(~input_layer[429]),
      .y(Y[1290]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1291_1
  function_186 neuron1291_1 (
      .a(input_layer[1312]),
      .b(~input_layer[362]),
      .c(input_layer[487]),
      .d(~input_layer[1337]),
      .y(Y[1291]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1292_1
  function_4 neuron1292_1 (
      .a(~input_layer[423]),
      .b(~input_layer[1433]),
      .c(~input_layer[230]),
      .d(~input_layer[123]),
      .e(~input_layer[1208]),
      .y(Y[1292]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1293_1
  function_27 neuron1293_1 (
      .a(~input_layer[1194]),
      .b(~input_layer[197]),
      .c(~input_layer[389]),
      .y(Y[1293]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1294_1
  function_47 neuron1294_1 (
      .a(input_layer[309]),
      .b(input_layer[411]),
      .c(input_layer[664]),
      .d(input_layer[733]),
      .e(input_layer[1162]),
      .y(Y[1294]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1295_1
  function_172 neuron1295_1 (
      .a(~input_layer[807]),
      .b(~input_layer[609]),
      .c(~input_layer[1112]),
      .d(input_layer[1034]),
      .e(~input_layer[1080]),
      .f(~input_layer[1293]),
      .y(Y[1295]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1296_1
  function_42 neuron1296_1 (
      .a(input_layer[637]),
      .b(input_layer[689]),
      .c(input_layer[194]),
      .d(~input_layer[1090]),
      .y(Y[1296]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1297_1
  function_19 neuron1297_1 (
      .a(~input_layer[756]),
      .b(~input_layer[915]),
      .c(~input_layer[909]),
      .d(input_layer[395]),
      .y(Y[1297]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1298_1
  function_7 neuron1298_1 (
      .a(input_layer[869]),
      .b(~input_layer[879]),
      .c(input_layer[122]),
      .d(input_layer[988]),
      .y(Y[1298]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1299_1
  function_17 neuron1299_1 (
      .a(input_layer[1129]),
      .b(input_layer[1166]),
      .c(~input_layer[814]),
      .y(Y[1299]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1300_1
  function_29 neuron1300_1 (
      .a(~input_layer[1036]),
      .b(~input_layer[130]),
      .y(Y[1300]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1301_1
  function_3 neuron1301_1 (
      .a(~input_layer[551]),
      .b(~input_layer[522]),
      .c(~input_layer[1018]),
      .d(~input_layer[190]),
      .y(Y[1301]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1302_1
  function_299 neuron1302_1 (
      .a(~input_layer[868]),
      .b(~input_layer[1061]),
      .c(~input_layer[515]),
      .d(input_layer[886]),
      .e(input_layer[1026]),
      .y(Y[1302]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1303_1
  function_30 neuron1303_1 (
      .a(input_layer[246]),
      .b(input_layer[1165]),
      .c(input_layer[1164]),
      .d(~input_layer[1430]),
      .y(Y[1303]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1304_1
  function_46 neuron1304_1 (
      .a(input_layer[202]),
      .b(input_layer[813]),
      .c(input_layer[79]),
      .d(~input_layer[674]),
      .e(input_layer[503]),
      .y(Y[1304]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1305_1
  function_60 neuron1305_1 (
      .a(input_layer[721]),
      .b(~input_layer[383]),
      .c(input_layer[309]),
      .d(input_layer[79]),
      .e(input_layer[1477]),
      .y(Y[1305]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_362 for neuron1306_1
  function_362 neuron1306_1 (
      .a(input_layer[927]),
      .b(input_layer[462]),
      .c(~input_layer[686]),
      .d(~input_layer[1218]),
      .e(input_layer[1182]),
      .f(input_layer[840]),
      .y(Y[1306]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_173 for neuron1307_1
  function_173 neuron1307_1 (
      .a(~input_layer[192]),
      .b(~input_layer[151]),
      .c(input_layer[1372]),
      .d(input_layer[525]),
      .e(~input_layer[1043]),
      .y(Y[1307]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_338 for neuron1308_1
  function_338 neuron1308_1 (
      .a(input_layer[1283]),
      .b(~input_layer[957]),
      .c(~input_layer[877]),
      .d(input_layer[506]),
      .e(input_layer[1272]),
      .f(input_layer[1513]),
      .y(Y[1308]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1309_1
  function_48 neuron1309_1 (
      .a(input_layer[687]),
      .b(input_layer[583]),
      .c(input_layer[1474]),
      .d(~input_layer[1264]),
      .e(input_layer[219]),
      .y(Y[1309]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1310] = 1'b0;

  // instantiate function_37 for neuron1311_1
  function_37 neuron1311_1 (
      .a(input_layer[1089]),
      .b(input_layer[140]),
      .c(input_layer[196]),
      .d(input_layer[88]),
      .e(~input_layer[561]),
      .f(input_layer[760]),
      .y(Y[1311]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1312_1
  function_19 neuron1312_1 (
      .a(input_layer[592]),
      .b(~input_layer[1486]),
      .c(~input_layer[1531]),
      .d(~input_layer[822]),
      .y(Y[1312]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_363 for neuron1313_1
  function_363 neuron1313_1 (
      .a(~input_layer[636]),
      .b(~input_layer[888]),
      .c(~input_layer[972]),
      .d(input_layer[376]),
      .e(~input_layer[615]),
      .f(input_layer[367]),
      .y(Y[1313]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron1314_1
  function_119 neuron1314_1 (
      .a(input_layer[1152]),
      .b(~input_layer[1429]),
      .c(~input_layer[674]),
      .d(input_layer[1051]),
      .e(input_layer[1050]),
      .y(Y[1314]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_364 for neuron1315_1
  function_364 neuron1315_1 (
      .a(~input_layer[661]),
      .b(input_layer[1238]),
      .c(input_layer[239]),
      .d(input_layer[184]),
      .e(input_layer[3]),
      .f(input_layer[10]),
      .y(Y[1315]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_365 for neuron1316_1
  function_365 neuron1316_1 (
      .a(input_layer[376]),
      .b(~input_layer[1411]),
      .c(~input_layer[528]),
      .d(input_layer[1293]),
      .e(input_layer[1310]),
      .f(input_layer[763]),
      .y(Y[1316]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron1317_1
  function_202 neuron1317_1 (
      .a(~input_layer[1024]),
      .b(~input_layer[1128]),
      .c(input_layer[878]),
      .d(input_layer[764]),
      .e(~input_layer[631]),
      .f(input_layer[1552]),
      .y(Y[1317]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_285 for neuron1318_1
  function_285 neuron1318_1 (
      .a(~input_layer[660]),
      .b(input_layer[1138]),
      .c(~input_layer[986]),
      .d(~input_layer[1382]),
      .e(~input_layer[101]),
      .f(~input_layer[425]),
      .y(Y[1318]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_366 for neuron1319_1
  function_366 neuron1319_1 (
      .a(~input_layer[1159]),
      .b(input_layer[567]),
      .c(input_layer[708]),
      .d(input_layer[396]),
      .e(input_layer[525]),
      .f(input_layer[55]),
      .y(Y[1319]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1320_1
  function_60 neuron1320_1 (
      .a(input_layer[138]),
      .b(input_layer[1240]),
      .c(~input_layer[518]),
      .d(input_layer[348]),
      .e(~input_layer[1229]),
      .y(Y[1320]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron1321_1
  function_242 neuron1321_1 (
      .a(input_layer[244]),
      .b(input_layer[314]),
      .c(~input_layer[1333]),
      .d(input_layer[92]),
      .e(~input_layer[747]),
      .f(input_layer[624]),
      .y(Y[1321]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_367 for neuron1322_1
  function_367 neuron1322_1 (
      .a(input_layer[422]),
      .b(~input_layer[1100]),
      .c(~input_layer[1191]),
      .d(input_layer[781]),
      .e(~input_layer[906]),
      .f(input_layer[35]),
      .y(Y[1322]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1323_1
  function_55 neuron1323_1 (
      .a(~input_layer[541]),
      .b(~input_layer[197]),
      .c(input_layer[431]),
      .d(input_layer[467]),
      .e(input_layer[1318]),
      .y(Y[1323]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1324_1
  function_0 neuron1324_1 (
      .a(~input_layer[1048]),
      .b(~input_layer[890]),
      .c(~input_layer[370]),
      .d(~input_layer[1257]),
      .e(~input_layer[1260]),
      .y(Y[1324]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1325_1
  function_16 neuron1325_1 (
      .a(input_layer[854]),
      .b(~input_layer[922]),
      .y(Y[1325]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1326_1
  function_39 neuron1326_1 (
      .a(input_layer[1169]),
      .b(~input_layer[153]),
      .c(~input_layer[856]),
      .y(Y[1326]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_368 for neuron1327_1
  function_368 neuron1327_1 (
      .a(~input_layer[699]),
      .b(input_layer[1487]),
      .c(input_layer[1496]),
      .d(~input_layer[356]),
      .e(~input_layer[446]),
      .f(input_layer[1428]),
      .y(Y[1327]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_369 for neuron1328_1
  function_369 neuron1328_1 (
      .a(~input_layer[629]),
      .b(~input_layer[436]),
      .c(~input_layer[155]),
      .d(input_layer[294]),
      .e(input_layer[532]),
      .f(input_layer[233]),
      .y(Y[1328]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1329_1
  function_0 neuron1329_1 (
      .a(~input_layer[1299]),
      .b(~input_layer[534]),
      .c(~input_layer[1026]),
      .d(~input_layer[343]),
      .e(~input_layer[895]),
      .y(Y[1329]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron1330_1
  function_241 neuron1330_1 (
      .a(input_layer[764]),
      .b(input_layer[150]),
      .c(input_layer[1001]),
      .d(input_layer[1537]),
      .e(input_layer[1236]),
      .f(input_layer[1053]),
      .y(Y[1330]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_370 for neuron1331_1
  function_370 neuron1331_1 (
      .a(~input_layer[349]),
      .b(input_layer[824]),
      .c(input_layer[533]),
      .d(~input_layer[1139]),
      .e(~input_layer[462]),
      .f(input_layer[941]),
      .y(Y[1331]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1332_1
  function_12 neuron1332_1 (
      .a(~input_layer[1137]),
      .b(input_layer[399]),
      .c(input_layer[791]),
      .y(Y[1332]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_212 for neuron1333_1
  function_212 neuron1333_1 (
      .a(~input_layer[686]),
      .b(input_layer[241]),
      .c(input_layer[1333]),
      .d(input_layer[1294]),
      .e(~input_layer[90]),
      .y(Y[1333]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1334_1
  function_35 neuron1334_1 (
      .a(~input_layer[1110]),
      .b(~input_layer[820]),
      .c(~input_layer[891]),
      .d(input_layer[1247]),
      .e(~input_layer[515]),
      .y(Y[1334]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1335] = 1'b0;

  // instantiate function_282 for neuron1336_1
  function_282 neuron1336_1 (
      .a(input_layer[851]),
      .b(~input_layer[501]),
      .c(~input_layer[1356]),
      .d(~input_layer[628]),
      .e(input_layer[1338]),
      .f(~input_layer[409]),
      .y(Y[1336]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_371 for neuron1337_1
  function_371 neuron1337_1 (
      .a(~input_layer[318]),
      .b(input_layer[1482]),
      .c(~input_layer[677]),
      .d(input_layer[792]),
      .e(~input_layer[284]),
      .f(input_layer[1410]),
      .y(Y[1337]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_372 for neuron1338_1
  function_372 neuron1338_1 (
      .a(~input_layer[438]),
      .b(input_layer[204]),
      .c(input_layer[90]),
      .d(~input_layer[349]),
      .e(input_layer[74]),
      .f(~input_layer[564]),
      .y(Y[1338]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_373 for neuron1339_1
  function_373 neuron1339_1 (
      .a(input_layer[318]),
      .b(input_layer[1251]),
      .c(input_layer[675]),
      .d(~input_layer[684]),
      .e(~input_layer[742]),
      .f(~input_layer[102]),
      .y(Y[1339]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_374 for neuron1340_1
  function_374 neuron1340_1 (
      .a(~input_layer[1145]),
      .b(~input_layer[715]),
      .c(input_layer[421]),
      .d(~input_layer[450]),
      .e(input_layer[1061]),
      .f(~input_layer[968]),
      .y(Y[1340]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_375 for neuron1341_1
  function_375 neuron1341_1 (
      .a(input_layer[1438]),
      .b(~input_layer[643]),
      .c(~input_layer[1206]),
      .d(~input_layer[408]),
      .e(~input_layer[540]),
      .y(Y[1341]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1342_1
  function_149 neuron1342_1 (
      .a(input_layer[983]),
      .b(~input_layer[1198]),
      .c(~input_layer[91]),
      .d(input_layer[1536]),
      .y(Y[1342]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1343_1
  function_0 neuron1343_1 (
      .a(~input_layer[1277]),
      .b(~input_layer[857]),
      .c(~input_layer[216]),
      .d(input_layer[873]),
      .e(~input_layer[844]),
      .y(Y[1343]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1344_1
  function_42 neuron1344_1 (
      .a(input_layer[1482]),
      .b(input_layer[546]),
      .c(input_layer[747]),
      .d(input_layer[995]),
      .y(Y[1344]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_108 for neuron1345_1
  function_108 neuron1345_1 (
      .a(input_layer[347]),
      .b(~input_layer[1314]),
      .c(input_layer[919]),
      .d(input_layer[1111]),
      .e(input_layer[200]),
      .f(input_layer[1385]),
      .y(Y[1345]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1346] = 1'b1;

  // instantiate function_89 for neuron1347_1
  function_89 neuron1347_1 (
      .a(input_layer[1037]),
      .b(~input_layer[362]),
      .c(input_layer[593]),
      .d(~input_layer[948]),
      .e(~input_layer[684]),
      .y(Y[1347]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_206 for neuron1348_1
  function_206 neuron1348_1 (
      .a(~input_layer[144]),
      .b(~input_layer[1002]),
      .c(input_layer[1507]),
      .d(~input_layer[64]),
      .e(input_layer[59]),
      .f(input_layer[165]),
      .y(Y[1348]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1349_1
  function_26 neuron1349_1 (
      .a(~input_layer[831]),
      .y(Y[1349]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1350_1
  function_31 neuron1350_1 (
      .a(input_layer[1113]),
      .b(~input_layer[1544]),
      .c(~input_layer[620]),
      .d(~input_layer[533]),
      .y(Y[1350]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1351_1
  function_27 neuron1351_1 (
      .a(~input_layer[862]),
      .b(~input_layer[188]),
      .c(input_layer[532]),
      .y(Y[1351]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_376 for neuron1352_1
  function_376 neuron1352_1 (
      .a(~input_layer[888]),
      .b(~input_layer[969]),
      .c(input_layer[588]),
      .d(input_layer[1545]),
      .e(~input_layer[1189]),
      .f(input_layer[1551]),
      .y(Y[1352]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1353_1
  function_92 neuron1353_1 (
      .a(input_layer[320]),
      .b(input_layer[941]),
      .c(input_layer[888]),
      .d(input_layer[945]),
      .e(input_layer[1318]),
      .f(input_layer[1103]),
      .y(Y[1353]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_200 for neuron1354_1
  function_200 neuron1354_1 (
      .a(input_layer[1420]),
      .b(~input_layer[990]),
      .c(~input_layer[152]),
      .d(~input_layer[286]),
      .e(input_layer[660]),
      .f(~input_layer[1393]),
      .y(Y[1354]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1355_1
  function_39 neuron1355_1 (
      .a(~input_layer[997]),
      .b(input_layer[386]),
      .c(~input_layer[1500]),
      .y(Y[1355]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1356_1
  function_17 neuron1356_1 (
      .a(input_layer[821]),
      .b(~input_layer[552]),
      .c(input_layer[779]),
      .y(Y[1356]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1357_1
  function_44 neuron1357_1 (
      .a(~input_layer[210]),
      .b(input_layer[484]),
      .c(input_layer[376]),
      .d(input_layer[981]),
      .e(input_layer[954]),
      .y(Y[1357]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1358_1
  function_35 neuron1358_1 (
      .a(input_layer[748]),
      .b(~input_layer[129]),
      .c(~input_layer[1199]),
      .d(~input_layer[681]),
      .e(~input_layer[1095]),
      .y(Y[1358]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1359_1
  function_20 neuron1359_1 (
      .a(~input_layer[647]),
      .b(~input_layer[438]),
      .c(~input_layer[1393]),
      .d(input_layer[908]),
      .e(input_layer[1092]),
      .y(Y[1359]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron1360_1
  function_36 neuron1360_1 (
      .a(input_layer[1185]),
      .b(input_layer[358]),
      .c(input_layer[1239]),
      .d(~input_layer[868]),
      .e(input_layer[254]),
      .f(~input_layer[23]),
      .y(Y[1360]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1361_1
  function_29 neuron1361_1 (
      .a(~input_layer[816]),
      .b(~input_layer[1419]),
      .y(Y[1361]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1362_1
  function_214 neuron1362_1 (
      .a(input_layer[137]),
      .b(~input_layer[696]),
      .c(input_layer[857]),
      .d(input_layer[1392]),
      .e(input_layer[1360]),
      .f(input_layer[338]),
      .y(Y[1362]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1363_1
  function_60 neuron1363_1 (
      .a(input_layer[858]),
      .b(input_layer[923]),
      .c(input_layer[1220]),
      .d(~input_layer[1409]),
      .e(input_layer[98]),
      .y(Y[1363]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1364_1
  function_19 neuron1364_1 (
      .a(~input_layer[298]),
      .b(~input_layer[921]),
      .c(~input_layer[1326]),
      .d(~input_layer[1264]),
      .y(Y[1364]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1365_1
  function_48 neuron1365_1 (
      .a(input_layer[549]),
      .b(input_layer[942]),
      .c(input_layer[724]),
      .d(input_layer[768]),
      .e(~input_layer[901]),
      .y(Y[1365]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron1366_1
  function_155 neuron1366_1 (
      .a(~input_layer[406]),
      .b(~input_layer[653]),
      .c(~input_layer[569]),
      .d(~input_layer[847]),
      .e(~input_layer[1553]),
      .f(~input_layer[163]),
      .y(Y[1366]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1367_1
  function_26 neuron1367_1 (
      .a(input_layer[757]),
      .y(Y[1367]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1368_1
  function_78 neuron1368_1 (
      .a(~input_layer[883]),
      .b(input_layer[311]),
      .c(~input_layer[881]),
      .d(~input_layer[620]),
      .e(~input_layer[1174]),
      .f(~input_layer[953]),
      .y(Y[1368]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1369_1
  function_167 neuron1369_1 (
      .a(input_layer[1136]),
      .b(input_layer[1053]),
      .c(input_layer[1327]),
      .d(input_layer[321]),
      .e(~input_layer[1434]),
      .y(Y[1369]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1370_1
  function_29 neuron1370_1 (
      .a(~input_layer[1076]),
      .b(~input_layer[320]),
      .y(Y[1370]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1371_1
  function_28 neuron1371_1 (
      .a(~input_layer[464]),
      .b(~input_layer[526]),
      .c(~input_layer[1049]),
      .d(~input_layer[1055]),
      .e(~input_layer[1115]),
      .f(~input_layer[719]),
      .y(Y[1371]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_377 for neuron1372_1
  function_377 neuron1372_1 (
      .a(~input_layer[606]),
      .b(input_layer[1126]),
      .c(input_layer[1541]),
      .d(~input_layer[1210]),
      .e(input_layer[505]),
      .f(~input_layer[614]),
      .y(Y[1372]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_349 for neuron1373_1
  function_349 neuron1373_1 (
      .a(input_layer[275]),
      .b(input_layer[1469]),
      .c(~input_layer[1081]),
      .d(~input_layer[304]),
      .e(input_layer[519]),
      .y(Y[1373]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1374_1
  function_45 neuron1374_1 (
      .a(input_layer[550]),
      .b(input_layer[875]),
      .c(input_layer[918]),
      .d(~input_layer[700]),
      .e(input_layer[659]),
      .f(~input_layer[1194]),
      .y(Y[1374]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1375_1
  function_27 neuron1375_1 (
      .a(input_layer[522]),
      .b(~input_layer[977]),
      .c(~input_layer[1162]),
      .y(Y[1375]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1376_1
  function_7 neuron1376_1 (
      .a(~input_layer[929]),
      .b(input_layer[1544]),
      .c(input_layer[1225]),
      .d(~input_layer[734]),
      .y(Y[1376]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1377_1
  function_97 neuron1377_1 (
      .a(input_layer[1436]),
      .b(~input_layer[1015]),
      .c(~input_layer[1171]),
      .d(~input_layer[1227]),
      .e(~input_layer[990]),
      .y(Y[1377]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1378_1
  function_90 neuron1378_1 (
      .a(~input_layer[1310]),
      .b(~input_layer[414]),
      .c(~input_layer[605]),
      .d(input_layer[676]),
      .e(~input_layer[1285]),
      .y(Y[1378]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1379_1
  function_30 neuron1379_1 (
      .a(input_layer[1075]),
      .b(input_layer[1439]),
      .c(~input_layer[861]),
      .d(~input_layer[940]),
      .y(Y[1379]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_378 for neuron1380_1
  function_378 neuron1380_1 (
      .a(~input_layer[135]),
      .b(input_layer[958]),
      .c(~input_layer[184]),
      .d(input_layer[355]),
      .e(input_layer[1302]),
      .f(input_layer[709]),
      .y(Y[1380]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1381_1
  function_167 neuron1381_1 (
      .a(input_layer[319]),
      .b(input_layer[1051]),
      .c(input_layer[432]),
      .d(input_layer[593]),
      .e(~input_layer[375]),
      .y(Y[1381]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1382_1
  function_334 neuron1382_1 (
      .a(input_layer[924]),
      .b(~input_layer[1137]),
      .c(input_layer[178]),
      .d(input_layer[1063]),
      .e(input_layer[894]),
      .y(Y[1382]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron1383_1
  function_157 neuron1383_1 (
      .a(input_layer[924]),
      .b(~input_layer[656]),
      .c(~input_layer[744]),
      .d(~input_layer[596]),
      .e(input_layer[730]),
      .f(input_layer[673]),
      .y(Y[1383]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1384_1
  function_17 neuron1384_1 (
      .a(input_layer[477]),
      .b(input_layer[1536]),
      .c(input_layer[587]),
      .y(Y[1384]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_379 for neuron1385_1
  function_379 neuron1385_1 (
      .a(~input_layer[1317]),
      .b(~input_layer[1372]),
      .c(input_layer[817]),
      .d(~input_layer[465]),
      .e(~input_layer[410]),
      .f(input_layer[651]),
      .y(Y[1385]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1386_1
  function_78 neuron1386_1 (
      .a(~input_layer[1365]),
      .b(~input_layer[549]),
      .c(input_layer[870]),
      .d(~input_layer[736]),
      .e(~input_layer[1063]),
      .f(~input_layer[950]),
      .y(Y[1386]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1387_1
  function_16 neuron1387_1 (
      .a(input_layer[857]),
      .b(input_layer[1443]),
      .y(Y[1387]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1388_1
  function_146 neuron1388_1 (
      .a(input_layer[1374]),
      .b(input_layer[1308]),
      .c(input_layer[444]),
      .d(~input_layer[716]),
      .e(input_layer[346]),
      .f(input_layer[733]),
      .y(Y[1388]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1389_1
  function_12 neuron1389_1 (
      .a(input_layer[864]),
      .b(~input_layer[767]),
      .c(input_layer[500]),
      .y(Y[1389]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron1390_1
  function_93 neuron1390_1 (
      .a(~input_layer[974]),
      .b(input_layer[399]),
      .c(input_layer[193]),
      .d(input_layer[1247]),
      .e(~input_layer[163]),
      .y(Y[1390]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1391_1
  function_19 neuron1391_1 (
      .a(~input_layer[934]),
      .b(~input_layer[1048]),
      .c(input_layer[754]),
      .d(~input_layer[1498]),
      .y(Y[1391]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_313 for neuron1392_1
  function_313 neuron1392_1 (
      .a(~input_layer[1435]),
      .b(input_layer[1100]),
      .c(input_layer[81]),
      .d(input_layer[618]),
      .e(~input_layer[586]),
      .f(~input_layer[1462]),
      .y(Y[1392]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_295 for neuron1393_1
  function_295 neuron1393_1 (
      .a(~input_layer[715]),
      .b(~input_layer[1055]),
      .c(input_layer[385]),
      .d(input_layer[328]),
      .e(input_layer[1371]),
      .f(input_layer[791]),
      .y(Y[1393]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1394_1
  function_3 neuron1394_1 (
      .a(~input_layer[1018]),
      .b(~input_layer[762]),
      .c(~input_layer[297]),
      .d(~input_layer[1165]),
      .y(Y[1394]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron1395_1
  function_152 neuron1395_1 (
      .a(~input_layer[1039]),
      .b(~input_layer[192]),
      .c(~input_layer[1165]),
      .d(input_layer[287]),
      .e(~input_layer[1014]),
      .y(Y[1395]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1396_1
  function_149 neuron1396_1 (
      .a(~input_layer[1276]),
      .b(~input_layer[746]),
      .c(~input_layer[331]),
      .d(input_layer[1545]),
      .y(Y[1396]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1397_1
  function_16 neuron1397_1 (
      .a(input_layer[974]),
      .b(input_layer[1333]),
      .y(Y[1397]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_380 for neuron1398_1
  function_380 neuron1398_1 (
      .a(input_layer[1159]),
      .b(~input_layer[470]),
      .c(~input_layer[1413]),
      .d(~input_layer[1226]),
      .e(input_layer[869]),
      .f(input_layer[179]),
      .y(Y[1398]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1399_1
  function_42 neuron1399_1 (
      .a(input_layer[883]),
      .b(input_layer[445]),
      .c(input_layer[1048]),
      .d(input_layer[1003]),
      .y(Y[1399]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1400_1
  function_17 neuron1400_1 (
      .a(input_layer[130]),
      .b(input_layer[703]),
      .c(input_layer[1474]),
      .y(Y[1400]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1401_1
  function_17 neuron1401_1 (
      .a(input_layer[184]),
      .b(input_layer[1124]),
      .c(~input_layer[430]),
      .y(Y[1401]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1402_1
  function_67 neuron1402_1 (
      .a(~input_layer[1359]),
      .b(~input_layer[1418]),
      .c(~input_layer[1248]),
      .d(input_layer[1206]),
      .e(~input_layer[289]),
      .y(Y[1402]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_238 for neuron1403_1
  function_238 neuron1403_1 (
      .a(input_layer[717]),
      .b(~input_layer[1224]),
      .c(~input_layer[1155]),
      .d(input_layer[1532]),
      .e(input_layer[215]),
      .y(Y[1403]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1404_1
  function_35 neuron1404_1 (
      .a(~input_layer[1075]),
      .b(input_layer[864]),
      .c(~input_layer[566]),
      .d(~input_layer[235]),
      .e(~input_layer[702]),
      .y(Y[1404]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron1405_1
  function_221 neuron1405_1 (
      .a(input_layer[312]),
      .b(input_layer[609]),
      .c(input_layer[265]),
      .d(~input_layer[1224]),
      .e(input_layer[513]),
      .f(~input_layer[1273]),
      .y(Y[1405]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1406_1
  function_60 neuron1406_1 (
      .a(input_layer[207]),
      .b(~input_layer[918]),
      .c(input_layer[441]),
      .d(~input_layer[976]),
      .e(input_layer[960]),
      .y(Y[1406]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1407_1
  function_31 neuron1407_1 (
      .a(~input_layer[1191]),
      .b(~input_layer[237]),
      .c(input_layer[681]),
      .d(input_layer[565]),
      .y(Y[1407]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1408_1
  function_146 neuron1408_1 (
      .a(input_layer[1485]),
      .b(input_layer[1191]),
      .c(input_layer[445]),
      .d(input_layer[565]),
      .e(~input_layer[379]),
      .f(input_layer[563]),
      .y(Y[1408]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_381 for neuron1409_1
  function_381 neuron1409_1 (
      .a(~input_layer[577]),
      .b(~input_layer[1441]),
      .c(input_layer[1107]),
      .d(input_layer[255]),
      .e(input_layer[1020]),
      .f(~input_layer[564]),
      .y(Y[1409]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1410_1
  function_181 neuron1410_1 (
      .a(input_layer[631]),
      .b(input_layer[680]),
      .c(~input_layer[1280]),
      .d(input_layer[1406]),
      .e(~input_layer[1412]),
      .y(Y[1410]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1411_1
  function_24 neuron1411_1 (
      .a(~input_layer[801]),
      .b(input_layer[1359]),
      .c(~input_layer[1385]),
      .y(Y[1411]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1412_1
  function_27 neuron1412_1 (
      .a(~input_layer[1430]),
      .b(input_layer[1146]),
      .c(~input_layer[492]),
      .y(Y[1412]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1413_1
  function_42 neuron1413_1 (
      .a(input_layer[832]),
      .b(input_layer[344]),
      .c(input_layer[233]),
      .d(input_layer[179]),
      .y(Y[1413]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron1414_1
  function_82 neuron1414_1 (
      .a(~input_layer[795]),
      .b(input_layer[350]),
      .c(input_layer[1263]),
      .d(~input_layer[587]),
      .e(~input_layer[620]),
      .f(~input_layer[1008]),
      .y(Y[1414]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1415_1
  function_17 neuron1415_1 (
      .a(~input_layer[908]),
      .b(input_layer[781]),
      .c(input_layer[1466]),
      .y(Y[1415]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1416_1
  function_12 neuron1416_1 (
      .a(input_layer[1083]),
      .b(~input_layer[916]),
      .c(input_layer[571]),
      .y(Y[1416]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1417_1
  function_55 neuron1417_1 (
      .a(~input_layer[553]),
      .b(input_layer[1142]),
      .c(~input_layer[1441]),
      .d(~input_layer[795]),
      .e(~input_layer[1443]),
      .y(Y[1417]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1418_1
  function_0 neuron1418_1 (
      .a(~input_layer[434]),
      .b(input_layer[588]),
      .c(~input_layer[1430]),
      .d(~input_layer[1138]),
      .e(~input_layer[124]),
      .y(Y[1418]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1419_1
  function_29 neuron1419_1 (
      .a(~input_layer[154]),
      .b(~input_layer[80]),
      .y(Y[1419]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron1420_1
  function_74 neuron1420_1 (
      .a(~input_layer[1278]),
      .b(~input_layer[182]),
      .c(~input_layer[481]),
      .d(~input_layer[466]),
      .e(~input_layer[230]),
      .f(input_layer[1232]),
      .y(Y[1420]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1421_1
  function_26 neuron1421_1 (
      .a(input_layer[749]),
      .y(Y[1421]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1422_1
  function_214 neuron1422_1 (
      .a(input_layer[851]),
      .b(input_layer[715]),
      .c(input_layer[322]),
      .d(~input_layer[1522]),
      .e(input_layer[157]),
      .f(~input_layer[449]),
      .y(Y[1422]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1423_1
  function_90 neuron1423_1 (
      .a(~input_layer[1149]),
      .b(~input_layer[1070]),
      .c(~input_layer[255]),
      .d(~input_layer[373]),
      .e(~input_layer[1306]),
      .y(Y[1423]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1424_1
  function_106 neuron1424_1 (
      .a(~input_layer[310]),
      .b(input_layer[1259]),
      .c(input_layer[1535]),
      .d(~input_layer[299]),
      .y(Y[1424]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1425_1
  function_172 neuron1425_1 (
      .a(~input_layer[467]),
      .b(~input_layer[1105]),
      .c(~input_layer[1185]),
      .d(~input_layer[253]),
      .e(~input_layer[1173]),
      .f(input_layer[1313]),
      .y(Y[1425]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1426_1
  function_3 neuron1426_1 (
      .a(~input_layer[1250]),
      .b(~input_layer[209]),
      .c(~input_layer[345]),
      .d(~input_layer[780]),
      .y(Y[1426]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1427_1
  function_319 neuron1427_1 (
      .a(input_layer[1489]),
      .b(input_layer[650]),
      .c(~input_layer[200]),
      .d(~input_layer[632]),
      .e(input_layer[1372]),
      .f(input_layer[287]),
      .y(Y[1427]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1428_1
  function_11 neuron1428_1 (
      .a(~input_layer[496]),
      .b(~input_layer[1358]),
      .c(input_layer[1442]),
      .d(~input_layer[1467]),
      .y(Y[1428]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1429_1
  function_67 neuron1429_1 (
      .a(~input_layer[469]),
      .b(~input_layer[214]),
      .c(~input_layer[711]),
      .d(~input_layer[937]),
      .e(~input_layer[402]),
      .y(Y[1429]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron1430_1
  function_119 neuron1430_1 (
      .a(~input_layer[743]),
      .b(~input_layer[1315]),
      .c(input_layer[563]),
      .d(~input_layer[1389]),
      .e(~input_layer[1404]),
      .y(Y[1430]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1431_1
  function_126 neuron1431_1 (
      .a(~input_layer[445]),
      .b(input_layer[905]),
      .c(~input_layer[551]),
      .d(~input_layer[1466]),
      .e(~input_layer[1292]),
      .y(Y[1431]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_382 for neuron1432_1
  function_382 neuron1432_1 (
      .a(~input_layer[1113]),
      .b(~input_layer[469]),
      .c(~input_layer[1196]),
      .d(~input_layer[253]),
      .e(~input_layer[352]),
      .f(~input_layer[222]),
      .y(Y[1432]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1433_1
  function_24 neuron1433_1 (
      .a(input_layer[750]),
      .b(~input_layer[259]),
      .c(input_layer[578]),
      .y(Y[1433]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_218 for neuron1434_1
  function_218 neuron1434_1 (
      .a(input_layer[1115]),
      .b(~input_layer[588]),
      .c(input_layer[1117]),
      .d(~input_layer[1068]),
      .e(~input_layer[444]),
      .y(Y[1434]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1435_1
  function_148 neuron1435_1 (
      .a(input_layer[496]),
      .b(input_layer[904]),
      .c(~input_layer[662]),
      .d(~input_layer[1444]),
      .e(~input_layer[24]),
      .f(~input_layer[1567]),
      .y(Y[1435]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_383 for neuron1436_1
  function_383 neuron1436_1 (
      .a(~input_layer[712]),
      .b(input_layer[927]),
      .c(input_layer[501]),
      .d(~input_layer[629]),
      .e(~input_layer[736]),
      .f(~input_layer[1402]),
      .y(Y[1436]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1437_1
  function_167 neuron1437_1 (
      .a(input_layer[352]),
      .b(input_layer[252]),
      .c(input_layer[1237]),
      .d(~input_layer[582]),
      .e(~input_layer[876]),
      .y(Y[1437]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1438_1
  function_39 neuron1438_1 (
      .a(input_layer[440]),
      .b(~input_layer[350]),
      .c(input_layer[1323]),
      .y(Y[1438]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1439_1
  function_26 neuron1439_1 (
      .a(~input_layer[423]),
      .y(Y[1439]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1440_1
  function_17 neuron1440_1 (
      .a(input_layer[146]),
      .b(input_layer[889]),
      .c(~input_layer[412]),
      .y(Y[1440]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron1441_1
  function_165 neuron1441_1 (
      .a(~input_layer[998]),
      .b(~input_layer[1219]),
      .c(input_layer[623]),
      .d(input_layer[1247]),
      .e(~input_layer[21]),
      .y(Y[1441]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_384 for neuron1442_1
  function_384 neuron1442_1 (
      .a(input_layer[1057]),
      .b(input_layer[920]),
      .c(~input_layer[397]),
      .d(~input_layer[816]),
      .e(~input_layer[988]),
      .f(~input_layer[521]),
      .y(Y[1442]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1443_1
  function_16 neuron1443_1 (
      .a(input_layer[529]),
      .b(input_layer[945]),
      .y(Y[1443]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_385 for neuron1444_1
  function_385 neuron1444_1 (
      .a(input_layer[1143]),
      .b(input_layer[1195]),
      .c(~input_layer[1374]),
      .d(~input_layer[516]),
      .e(input_layer[1392]),
      .f(~input_layer[139]),
      .y(Y[1444]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1445_1
  function_149 neuron1445_1 (
      .a(input_layer[1198]),
      .b(~input_layer[1529]),
      .c(input_layer[918]),
      .d(~input_layer[1114]),
      .y(Y[1445]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1446_1
  function_16 neuron1446_1 (
      .a(~input_layer[1036]),
      .b(input_layer[1016]),
      .y(Y[1446]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_386 for neuron1447_1
  function_386 neuron1447_1 (
      .a(input_layer[1055]),
      .b(~input_layer[155]),
      .c(input_layer[302]),
      .d(~input_layer[510]),
      .e(input_layer[196]),
      .f(input_layer[951]),
      .y(Y[1447]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_387 for neuron1448_1
  function_387 neuron1448_1 (
      .a(input_layer[694]),
      .b(~input_layer[765]),
      .c(~input_layer[1413]),
      .d(input_layer[753]),
      .e(~input_layer[1359]),
      .f(input_layer[433]),
      .y(Y[1448]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1449_1
  function_214 neuron1449_1 (
      .a(input_layer[608]),
      .b(input_layer[1438]),
      .c(input_layer[1362]),
      .d(~input_layer[1329]),
      .e(~input_layer[271]),
      .f(input_layer[759]),
      .y(Y[1449]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_238 for neuron1450_1
  function_238 neuron1450_1 (
      .a(input_layer[1091]),
      .b(input_layer[509]),
      .c(~input_layer[237]),
      .d(input_layer[333]),
      .e(~input_layer[317]),
      .y(Y[1450]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1451_1
  function_89 neuron1451_1 (
      .a(~input_layer[1217]),
      .b(input_layer[1546]),
      .c(input_layer[762]),
      .d(input_layer[1522]),
      .e(~input_layer[187]),
      .y(Y[1451]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1452_1
  function_148 neuron1452_1 (
      .a(input_layer[1415]),
      .b(~input_layer[756]),
      .c(input_layer[274]),
      .d(input_layer[1107]),
      .e(input_layer[1023]),
      .f(~input_layer[671]),
      .y(Y[1452]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_388 for neuron1453_1
  function_388 neuron1453_1 (
      .a(~input_layer[795]),
      .b(input_layer[1423]),
      .c(~input_layer[1034]),
      .d(input_layer[1421]),
      .e(input_layer[1196]),
      .f(input_layer[304]),
      .y(Y[1453]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_389 for neuron1454_1
  function_389 neuron1454_1 (
      .a(input_layer[1032]),
      .b(input_layer[1305]),
      .c(input_layer[431]),
      .d(~input_layer[343]),
      .e(input_layer[1219]),
      .f(input_layer[3]),
      .y(Y[1454]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1455_1
  function_48 neuron1455_1 (
      .a(input_layer[1136]),
      .b(input_layer[1143]),
      .c(input_layer[1535]),
      .d(input_layer[1104]),
      .e(~input_layer[824]),
      .y(Y[1455]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_367 for neuron1456_1
  function_367 neuron1456_1 (
      .a(input_layer[498]),
      .b(~input_layer[1538]),
      .c(~input_layer[128]),
      .d(~input_layer[95]),
      .e(~input_layer[345]),
      .f(input_layer[1179]),
      .y(Y[1456]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_390 for neuron1457_1
  function_390 neuron1457_1 (
      .a(input_layer[1247]),
      .b(~input_layer[142]),
      .c(~input_layer[137]),
      .d(input_layer[364]),
      .e(~input_layer[1148]),
      .f(~input_layer[1295]),
      .y(Y[1457]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_391 for neuron1458_1
  function_391 neuron1458_1 (
      .a(input_layer[693]),
      .b(~input_layer[1237]),
      .c(~input_layer[1317]),
      .d(~input_layer[1004]),
      .e(~input_layer[606]),
      .f(~input_layer[467]),
      .y(Y[1458]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron1459_1
  function_119 neuron1459_1 (
      .a(~input_layer[808]),
      .b(~input_layer[979]),
      .c(input_layer[1483]),
      .d(input_layer[1550]),
      .e(input_layer[637]),
      .y(Y[1459]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_383 for neuron1460_1
  function_383 neuron1460_1 (
      .a(input_layer[749]),
      .b(~input_layer[1279]),
      .c(~input_layer[1029]),
      .d(input_layer[826]),
      .e(~input_layer[248]),
      .f(input_layer[184]),
      .y(Y[1460]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1461_1
  function_29 neuron1461_1 (
      .a(input_layer[799]),
      .b(~input_layer[958]),
      .y(Y[1461]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1462_1
  function_169 neuron1462_1 (
      .a(~input_layer[1130]),
      .b(input_layer[1030]),
      .c(~input_layer[1156]),
      .d(~input_layer[363]),
      .e(~input_layer[847]),
      .f(~input_layer[503]),
      .y(Y[1462]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron1463_1
  function_36 neuron1463_1 (
      .a(input_layer[204]),
      .b(input_layer[238]),
      .c(input_layer[890]),
      .d(input_layer[1012]),
      .e(~input_layer[809]),
      .f(~input_layer[1423]),
      .y(Y[1463]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1464_1
  function_12 neuron1464_1 (
      .a(~input_layer[424]),
      .b(input_layer[852]),
      .c(input_layer[884]),
      .y(Y[1464]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1465_1
  function_47 neuron1465_1 (
      .a(input_layer[967]),
      .b(input_layer[834]),
      .c(input_layer[467]),
      .d(input_layer[1236]),
      .e(input_layer[988]),
      .y(Y[1465]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_23 for neuron1466_1
  function_23 neuron1466_1 (
      .a(input_layer[1368]),
      .b(~input_layer[131]),
      .c(input_layer[791]),
      .d(input_layer[955]),
      .e(~input_layer[1257]),
      .f(input_layer[896]),
      .y(Y[1466]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_235 for neuron1467_1
  function_235 neuron1467_1 (
      .a(~input_layer[630]),
      .b(~input_layer[805]),
      .c(input_layer[353]),
      .d(~input_layer[273]),
      .e(input_layer[1489]),
      .y(Y[1467]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1468_1
  function_0 neuron1468_1 (
      .a(~input_layer[1239]),
      .b(input_layer[1142]),
      .c(~input_layer[1192]),
      .d(~input_layer[1218]),
      .e(~input_layer[1498]),
      .y(Y[1468]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1469_1
  function_67 neuron1469_1 (
      .a(~input_layer[152]),
      .b(~input_layer[130]),
      .c(~input_layer[1445]),
      .d(~input_layer[389]),
      .e(~input_layer[233]),
      .y(Y[1469]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1470_1
  function_95 neuron1470_1 (
      .a(~input_layer[1167]),
      .b(input_layer[665]),
      .c(input_layer[1434]),
      .d(~input_layer[722]),
      .y(Y[1470]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron1471_1
  function_157 neuron1471_1 (
      .a(input_layer[314]),
      .b(~input_layer[1281]),
      .c(input_layer[1020]),
      .d(input_layer[1303]),
      .e(input_layer[900]),
      .f(~input_layer[1464]),
      .y(Y[1471]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_392 for neuron1472_1
  function_392 neuron1472_1 (
      .a(~input_layer[939]),
      .b(~input_layer[138]),
      .c(input_layer[708]),
      .d(~input_layer[732]),
      .e(input_layer[1391]),
      .f(input_layer[653]),
      .y(Y[1472]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1473_1
  function_92 neuron1473_1 (
      .a(input_layer[540]),
      .b(input_layer[497]),
      .c(input_layer[603]),
      .d(input_layer[949]),
      .e(~input_layer[1208]),
      .f(~input_layer[743]),
      .y(Y[1473]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1474_1
  function_12 neuron1474_1 (
      .a(input_layer[818]),
      .b(~input_layer[661]),
      .c(~input_layer[713]),
      .y(Y[1474]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1475_1
  function_27 neuron1475_1 (
      .a(~input_layer[307]),
      .b(input_layer[480]),
      .c(~input_layer[1027]),
      .y(Y[1475]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1476_1
  function_186 neuron1476_1 (
      .a(input_layer[602]),
      .b(input_layer[971]),
      .c(~input_layer[1535]),
      .d(~input_layer[1180]),
      .y(Y[1476]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_393 for neuron1477_1
  function_393 neuron1477_1 (
      .a(input_layer[553]),
      .b(~input_layer[1301]),
      .c(~input_layer[475]),
      .d(~input_layer[303]),
      .e(~input_layer[678]),
      .f(input_layer[963]),
      .y(Y[1477]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1478_1
  function_26 neuron1478_1 (
      .a(~input_layer[1323]),
      .y(Y[1478]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1479_1
  function_29 neuron1479_1 (
      .a(input_layer[969]),
      .b(~input_layer[567]),
      .y(Y[1479]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1480_1
  function_95 neuron1480_1 (
      .a(~input_layer[591]),
      .b(input_layer[547]),
      .c(~input_layer[195]),
      .d(input_layer[929]),
      .y(Y[1480]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1481_1
  function_39 neuron1481_1 (
      .a(input_layer[299]),
      .b(input_layer[638]),
      .c(~input_layer[565]),
      .y(Y[1481]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_305 for neuron1482_1
  function_305 neuron1482_1 (
      .a(input_layer[660]),
      .b(~input_layer[1192]),
      .c(~input_layer[268]),
      .d(~input_layer[332]),
      .e(input_layer[619]),
      .y(Y[1482]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1483_1
  function_46 neuron1483_1 (
      .a(input_layer[516]),
      .b(input_layer[465]),
      .c(input_layer[1029]),
      .d(~input_layer[1237]),
      .e(input_layer[672]),
      .y(Y[1483]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron1484_1
  function_70 neuron1484_1 (
      .a(~input_layer[1243]),
      .b(input_layer[472]),
      .c(~input_layer[1257]),
      .d(~input_layer[908]),
      .e(input_layer[688]),
      .f(~input_layer[771]),
      .y(Y[1484]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1485_1
  function_42 neuron1485_1 (
      .a(input_layer[847]),
      .b(input_layer[347]),
      .c(~input_layer[756]),
      .d(~input_layer[1262]),
      .y(Y[1485]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1486_1
  function_299 neuron1486_1 (
      .a(~input_layer[416]),
      .b(~input_layer[1469]),
      .c(input_layer[461]),
      .d(~input_layer[600]),
      .e(~input_layer[712]),
      .y(Y[1486]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1487_1
  function_12 neuron1487_1 (
      .a(input_layer[1335]),
      .b(~input_layer[314]),
      .c(~input_layer[905]),
      .y(Y[1487]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_394 for neuron1488_1
  function_394 neuron1488_1 (
      .a(~input_layer[143]),
      .b(input_layer[1325]),
      .c(input_layer[1039]),
      .d(~input_layer[696]),
      .e(input_layer[41]),
      .f(input_layer[728]),
      .y(Y[1488]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1489_1
  function_39 neuron1489_1 (
      .a(input_layer[267]),
      .b(~input_layer[1358]),
      .c(~input_layer[1255]),
      .y(Y[1489]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1490_1
  function_46 neuron1490_1 (
      .a(input_layer[522]),
      .b(input_layer[1530]),
      .c(~input_layer[995]),
      .d(~input_layer[986]),
      .e(input_layer[128]),
      .y(Y[1490]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1491_1
  function_47 neuron1491_1 (
      .a(input_layer[359]),
      .b(input_layer[990]),
      .c(input_layer[467]),
      .d(input_layer[150]),
      .e(input_layer[1170]),
      .y(Y[1491]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1492_1
  function_42 neuron1492_1 (
      .a(input_layer[700]),
      .b(~input_layer[1312]),
      .c(input_layer[1180]),
      .d(input_layer[348]),
      .y(Y[1492]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_395 for neuron1493_1
  function_395 neuron1493_1 (
      .a(~input_layer[757]),
      .b(input_layer[986]),
      .c(~input_layer[626]),
      .d(input_layer[97]),
      .e(~input_layer[344]),
      .f(~input_layer[1340]),
      .y(Y[1493]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1494_1
  function_149 neuron1494_1 (
      .a(~input_layer[1079]),
      .b(~input_layer[208]),
      .c(input_layer[590]),
      .d(input_layer[1410]),
      .y(Y[1494]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1495_1
  function_8 neuron1495_1 (
      .a(input_layer[1493]),
      .b(~input_layer[1110]),
      .c(input_layer[1531]),
      .d(~input_layer[990]),
      .y(Y[1495]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1496_1
  function_12 neuron1496_1 (
      .a(~input_layer[813]),
      .b(input_layer[889]),
      .c(input_layer[890]),
      .y(Y[1496]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1497_1
  function_17 neuron1497_1 (
      .a(input_layer[598]),
      .b(input_layer[511]),
      .c(input_layer[1387]),
      .y(Y[1497]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1498_1
  function_35 neuron1498_1 (
      .a(~input_layer[977]),
      .b(~input_layer[500]),
      .c(~input_layer[829]),
      .d(input_layer[992]),
      .e(input_layer[1052]),
      .y(Y[1498]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1499_1
  function_27 neuron1499_1 (
      .a(~input_layer[257]),
      .b(~input_layer[311]),
      .c(~input_layer[757]),
      .y(Y[1499]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1500_1
  function_29 neuron1500_1 (
      .a(~input_layer[1127]),
      .b(input_layer[1248]),
      .y(Y[1500]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_302 for neuron1501_1
  function_302 neuron1501_1 (
      .a(~input_layer[538]),
      .b(input_layer[871]),
      .c(input_layer[692]),
      .d(~input_layer[988]),
      .e(~input_layer[232]),
      .f(input_layer[1493]),
      .y(Y[1501]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1502_1
  function_67 neuron1502_1 (
      .a(~input_layer[1115]),
      .b(~input_layer[242]),
      .c(~input_layer[265]),
      .d(input_layer[476]),
      .e(input_layer[762]),
      .y(Y[1502]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1503_1
  function_27 neuron1503_1 (
      .a(~input_layer[212]),
      .b(~input_layer[993]),
      .c(input_layer[598]),
      .y(Y[1503]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1504_1
  function_29 neuron1504_1 (
      .a(~input_layer[1193]),
      .b(input_layer[747]),
      .y(Y[1504]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1505_1
  function_146 neuron1505_1 (
      .a(input_layer[1483]),
      .b(input_layer[387]),
      .c(input_layer[1277]),
      .d(~input_layer[95]),
      .e(input_layer[789]),
      .f(~input_layer[630]),
      .y(Y[1505]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron1506_1
  function_234 neuron1506_1 (
      .a(input_layer[708]),
      .b(~input_layer[1164]),
      .c(~input_layer[1548]),
      .d(~input_layer[1258]),
      .e(~input_layer[295]),
      .f(input_layer[581]),
      .y(Y[1506]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1507_1
  function_16 neuron1507_1 (
      .a(~input_layer[1200]),
      .b(input_layer[848]),
      .y(Y[1507]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1508_1
  function_26 neuron1508_1 (
      .a(input_layer[712]),
      .y(Y[1508]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_338 for neuron1509_1
  function_338 neuron1509_1 (
      .a(input_layer[288]),
      .b(~input_layer[464]),
      .c(input_layer[772]),
      .d(input_layer[422]),
      .e(input_layer[1396]),
      .f(input_layer[1177]),
      .y(Y[1509]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1510_1
  function_39 neuron1510_1 (
      .a(~input_layer[1078]),
      .b(input_layer[1308]),
      .c(input_layer[520]),
      .y(Y[1510]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1511_1
  function_46 neuron1511_1 (
      .a(input_layer[555]),
      .b(input_layer[1186]),
      .c(input_layer[332]),
      .d(~input_layer[1497]),
      .e(input_layer[99]),
      .y(Y[1511]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_137 for neuron1512_1
  function_137 neuron1512_1 (
      .a(input_layer[199]),
      .b(input_layer[204]),
      .c(~input_layer[649]),
      .d(~input_layer[1112]),
      .e(input_layer[1095]),
      .y(Y[1512]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1513_1
  function_42 neuron1513_1 (
      .a(input_layer[767]),
      .b(input_layer[214]),
      .c(input_layer[1534]),
      .d(input_layer[288]),
      .y(Y[1513]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1514_1
  function_29 neuron1514_1 (
      .a(input_layer[193]),
      .b(~input_layer[1222]),
      .y(Y[1514]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1515_1
  function_330 neuron1515_1 (
      .a(~input_layer[1536]),
      .b(input_layer[210]),
      .c(~input_layer[651]),
      .d(~input_layer[874]),
      .e(~input_layer[52]),
      .y(Y[1515]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1516] = 1'b0;

  // instantiate function_91 for neuron1517_1
  function_91 neuron1517_1 (
      .a(input_layer[1256]),
      .b(~input_layer[1489]),
      .c(input_layer[696]),
      .d(input_layer[381]),
      .e(~input_layer[1392]),
      .y(Y[1517]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_396 for neuron1518_1
  function_396 neuron1518_1 (
      .a(input_layer[851]),
      .b(input_layer[601]),
      .c(input_layer[870]),
      .d(~input_layer[1189]),
      .e(~input_layer[779]),
      .y(Y[1518]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_397 for neuron1519_1
  function_397 neuron1519_1 (
      .a(~input_layer[1443]),
      .b(input_layer[889]),
      .c(input_layer[86]),
      .d(input_layer[71]),
      .e(~input_layer[500]),
      .y(Y[1519]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1520_1
  function_16 neuron1520_1 (
      .a(input_layer[1274]),
      .b(input_layer[1270]),
      .y(Y[1520]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron1521_1
  function_232 neuron1521_1 (
      .a(~input_layer[137]),
      .b(~input_layer[260]),
      .c(input_layer[1365]),
      .d(input_layer[628]),
      .e(input_layer[1266]),
      .f(~input_layer[65]),
      .y(Y[1521]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1522_1
  function_78 neuron1522_1 (
      .a(~input_layer[595]),
      .b(~input_layer[545]),
      .c(~input_layer[608]),
      .d(~input_layer[1421]),
      .e(~input_layer[911]),
      .f(input_layer[1119]),
      .y(Y[1522]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1523_1
  function_92 neuron1523_1 (
      .a(~input_layer[428]),
      .b(input_layer[1171]),
      .c(input_layer[1058]),
      .d(input_layer[89]),
      .e(~input_layer[368]),
      .f(input_layer[563]),
      .y(Y[1523]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1524_1
  function_12 neuron1524_1 (
      .a(~input_layer[743]),
      .b(input_layer[552]),
      .c(input_layer[435]),
      .y(Y[1524]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1525_1
  function_172 neuron1525_1 (
      .a(~input_layer[383]),
      .b(~input_layer[834]),
      .c(input_layer[706]),
      .d(~input_layer[89]),
      .e(~input_layer[619]),
      .f(~input_layer[826]),
      .y(Y[1525]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_217 for neuron1526_1
  function_217 neuron1526_1 (
      .a(input_layer[1083]),
      .b(input_layer[1036]),
      .c(~input_layer[805]),
      .d(~input_layer[543]),
      .e(input_layer[728]),
      .f(input_layer[47]),
      .y(Y[1526]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1527_1
  function_16 neuron1527_1 (
      .a(input_layer[692]),
      .b(input_layer[1393]),
      .y(Y[1527]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1528_1
  function_26 neuron1528_1 (
      .a(input_layer[1132]),
      .y(Y[1528]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron1529_1
  function_85 neuron1529_1 (
      .a(input_layer[481]),
      .b(input_layer[623]),
      .c(~input_layer[873]),
      .d(~input_layer[766]),
      .e(~input_layer[116]),
      .f(~input_layer[44]),
      .y(Y[1529]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1530_1
  function_12 neuron1530_1 (
      .a(input_layer[424]),
      .b(~input_layer[767]),
      .c(input_layer[836]),
      .y(Y[1530]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_177 for neuron1531_1
  function_177 neuron1531_1 (
      .a(~input_layer[715]),
      .b(input_layer[343]),
      .c(~input_layer[523]),
      .d(input_layer[556]),
      .e(input_layer[759]),
      .y(Y[1531]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1532_1
  function_26 neuron1532_1 (
      .a(input_layer[1373]),
      .y(Y[1532]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1533_1
  function_42 neuron1533_1 (
      .a(input_layer[188]),
      .b(input_layer[379]),
      .c(input_layer[1073]),
      .d(input_layer[1004]),
      .y(Y[1533]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1534_1
  function_31 neuron1534_1 (
      .a(~input_layer[327]),
      .b(input_layer[565]),
      .c(input_layer[888]),
      .d(~input_layer[124]),
      .y(Y[1534]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1535_1
  function_113 neuron1535_1 (
      .a(input_layer[1538]),
      .b(~input_layer[1036]),
      .c(input_layer[1447]),
      .d(~input_layer[1039]),
      .e(~input_layer[1334]),
      .y(Y[1535]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_22 for neuron1536_1
  function_22 neuron1536_1 (
      .a(input_layer[349]),
      .b(input_layer[1061]),
      .c(input_layer[450]),
      .d(~input_layer[1333]),
      .e(~input_layer[1448]),
      .f(input_layer[734]),
      .y(Y[1536]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1537_1
  function_3 neuron1537_1 (
      .a(~input_layer[1039]),
      .b(~input_layer[622]),
      .c(~input_layer[341]),
      .d(~input_layer[1007]),
      .y(Y[1537]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1538_1
  function_26 neuron1538_1 (
      .a(~input_layer[661]),
      .y(Y[1538]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_398 for neuron1539_1
  function_398 neuron1539_1 (
      .a(~input_layer[1196]),
      .b(input_layer[793]),
      .c(~input_layer[1161]),
      .d(~input_layer[1375]),
      .e(input_layer[369]),
      .f(~input_layer[210]),
      .y(Y[1539]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_368 for neuron1540_1
  function_368 neuron1540_1 (
      .a(input_layer[1113]),
      .b(input_layer[1473]),
      .c(~input_layer[212]),
      .d(input_layer[459]),
      .e(~input_layer[78]),
      .f(~input_layer[1306]),
      .y(Y[1540]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1541_1
  function_49 neuron1541_1 (
      .a(input_layer[757]),
      .b(~input_layer[1539]),
      .c(~input_layer[212]),
      .d(input_layer[1180]),
      .e(~input_layer[968]),
      .y(Y[1541]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_200 for neuron1542_1
  function_200 neuron1542_1 (
      .a(input_layer[746]),
      .b(~input_layer[1115]),
      .c(~input_layer[652]),
      .d(~input_layer[260]),
      .e(~input_layer[683]),
      .f(input_layer[431]),
      .y(Y[1542]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_399 for neuron1543_1
  function_399 neuron1543_1 (
      .a(~input_layer[811]),
      .b(input_layer[1151]),
      .c(input_layer[394]),
      .d(input_layer[344]),
      .e(input_layer[684]),
      .f(~input_layer[66]),
      .y(Y[1543]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_367 for neuron1544_1
  function_367 neuron1544_1 (
      .a(~input_layer[1073]),
      .b(~input_layer[757]),
      .c(~input_layer[1316]),
      .d(~input_layer[846]),
      .e(input_layer[1467]),
      .f(input_layer[1289]),
      .y(Y[1544]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1545_1
  function_47 neuron1545_1 (
      .a(input_layer[528]),
      .b(input_layer[519]),
      .c(input_layer[180]),
      .d(input_layer[1236]),
      .e(input_layer[459]),
      .y(Y[1545]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1546_1
  function_28 neuron1546_1 (
      .a(~input_layer[207]),
      .b(~input_layer[1298]),
      .c(~input_layer[1108]),
      .d(~input_layer[1147]),
      .e(~input_layer[1351]),
      .f(~input_layer[614]),
      .y(Y[1546]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron1547_1
  function_155 neuron1547_1 (
      .a(~input_layer[1139]),
      .b(~input_layer[1421]),
      .c(~input_layer[133]),
      .d(~input_layer[248]),
      .e(~input_layer[1047]),
      .f(input_layer[920]),
      .y(Y[1547]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1548_1
  function_3 neuron1548_1 (
      .a(~input_layer[187]),
      .b(~input_layer[935]),
      .c(input_layer[810]),
      .d(~input_layer[1350]),
      .y(Y[1548]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1549_1
  function_0 neuron1549_1 (
      .a(~input_layer[258]),
      .b(input_layer[421]),
      .c(~input_layer[155]),
      .d(~input_layer[957]),
      .e(~input_layer[1161]),
      .y(Y[1549]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1550_1
  function_48 neuron1550_1 (
      .a(input_layer[472]),
      .b(input_layer[585]),
      .c(input_layer[196]),
      .d(input_layer[1131]),
      .e(~input_layer[1304]),
      .y(Y[1550]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1551_1
  function_3 neuron1551_1 (
      .a(~input_layer[887]),
      .b(~input_layer[1297]),
      .c(~input_layer[180]),
      .d(~input_layer[1548]),
      .y(Y[1551]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1552_1
  function_307 neuron1552_1 (
      .a(~input_layer[908]),
      .b(input_layer[238]),
      .c(input_layer[1160]),
      .d(input_layer[780]),
      .e(input_layer[510]),
      .y(Y[1552]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1553_1
  function_146 neuron1553_1 (
      .a(input_layer[1480]),
      .b(input_layer[343]),
      .c(input_layer[1351]),
      .d(~input_layer[700]),
      .e(~input_layer[1219]),
      .f(input_layer[461]),
      .y(Y[1553]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1554_1
  function_12 neuron1554_1 (
      .a(~input_layer[368]),
      .b(input_layer[1532]),
      .c(input_layer[966]),
      .y(Y[1554]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1555_1
  function_11 neuron1555_1 (
      .a(~input_layer[768]),
      .b(~input_layer[246]),
      .c(input_layer[330]),
      .d(~input_layer[180]),
      .y(Y[1555]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1556_1
  function_16 neuron1556_1 (
      .a(input_layer[852]),
      .b(~input_layer[470]),
      .y(Y[1556]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1557_1
  function_28 neuron1557_1 (
      .a(~input_layer[299]),
      .b(~input_layer[1160]),
      .c(~input_layer[84]),
      .d(input_layer[880]),
      .e(~input_layer[78]),
      .f(~input_layer[360]),
      .y(Y[1557]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1558_1
  function_27 neuron1558_1 (
      .a(input_layer[698]),
      .b(~input_layer[1488]),
      .c(~input_layer[1416]),
      .y(Y[1558]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1559_1
  function_42 neuron1559_1 (
      .a(input_layer[251]),
      .b(input_layer[1360]),
      .c(input_layer[302]),
      .d(input_layer[1428]),
      .y(Y[1559]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1560_1
  function_186 neuron1560_1 (
      .a(input_layer[599]),
      .b(input_layer[459]),
      .c(~input_layer[1081]),
      .d(input_layer[819]),
      .y(Y[1560]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1561_1
  function_20 neuron1561_1 (
      .a(~input_layer[491]),
      .b(~input_layer[424]),
      .c(input_layer[657]),
      .d(input_layer[201]),
      .e(~input_layer[469]),
      .y(Y[1561]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_400 for neuron1562_1
  function_400 neuron1562_1 (
      .a(~input_layer[296]),
      .b(input_layer[1382]),
      .c(~input_layer[937]),
      .d(~input_layer[1181]),
      .e(~input_layer[97]),
      .f(input_layer[1413]),
      .y(Y[1562]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1563_1
  function_16 neuron1563_1 (
      .a(input_layer[682]),
      .b(~input_layer[308]),
      .y(Y[1563]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_255 for neuron1564_1
  function_255 neuron1564_1 (
      .a(input_layer[583]),
      .b(~input_layer[949]),
      .c(~input_layer[1046]),
      .d(~input_layer[291]),
      .e(input_layer[939]),
      .y(Y[1564]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1565_1
  function_42 neuron1565_1 (
      .a(input_layer[273]),
      .b(input_layer[189]),
      .c(~input_layer[817]),
      .d(input_layer[356]),
      .y(Y[1565]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_401 for neuron1566_1
  function_401 neuron1566_1 (
      .a(input_layer[910]),
      .b(~input_layer[629]),
      .c(input_layer[886]),
      .d(~input_layer[471]),
      .e(input_layer[248]),
      .f(~input_layer[615]),
      .y(Y[1566]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1567_1
  function_126 neuron1567_1 (
      .a(~input_layer[196]),
      .b(input_layer[850]),
      .c(~input_layer[1411]),
      .d(~input_layer[81]),
      .e(input_layer[384]),
      .y(Y[1567]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1568_1
  function_17 neuron1568_1 (
      .a(input_layer[211]),
      .b(input_layer[195]),
      .c(~input_layer[1214]),
      .y(Y[1568]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_383 for neuron1569_1
  function_383 neuron1569_1 (
      .a(~input_layer[1135]),
      .b(input_layer[1171]),
      .c(~input_layer[416]),
      .d(~input_layer[1374]),
      .e(input_layer[229]),
      .f(~input_layer[111]),
      .y(Y[1569]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_201 for neuron1570_1
  function_201 neuron1570_1 (
      .a(~input_layer[265]),
      .b(~input_layer[132]),
      .c(input_layer[1475]),
      .d(input_layer[403]),
      .e(~input_layer[256]),
      .f(~input_layer[64]),
      .y(Y[1570]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_402 for neuron1571_1
  function_402 neuron1571_1 (
      .a(input_layer[752]),
      .b(~input_layer[159]),
      .c(input_layer[343]),
      .d(input_layer[987]),
      .e(~input_layer[490]),
      .f(input_layer[994]),
      .y(Y[1571]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1572_1
  function_3 neuron1572_1 (
      .a(~input_layer[803]),
      .b(~input_layer[443]),
      .c(~input_layer[1298]),
      .d(input_layer[631]),
      .y(Y[1572]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_403 for neuron1573_1
  function_403 neuron1573_1 (
      .a(input_layer[767]),
      .b(~input_layer[436]),
      .c(~input_layer[1033]),
      .d(input_layer[1308]),
      .e(input_layer[468]),
      .f(~input_layer[1179]),
      .y(Y[1573]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron1574_1
  function_112 neuron1574_1 (
      .a(~input_layer[1305]),
      .b(~input_layer[575]),
      .c(~input_layer[285]),
      .d(input_layer[274]),
      .e(input_layer[1008]),
      .f(~input_layer[1520]),
      .y(Y[1574]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_404 for neuron1575_1
  function_404 neuron1575_1 (
      .a(input_layer[311]),
      .b(~input_layer[1545]),
      .c(~input_layer[94]),
      .d(input_layer[1145]),
      .e(~input_layer[1257]),
      .f(~input_layer[1064]),
      .y(Y[1575]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1576_1
  function_8 neuron1576_1 (
      .a(input_layer[793]),
      .b(~input_layer[1143]),
      .c(input_layer[1547]),
      .d(input_layer[946]),
      .y(Y[1576]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron1577_1
  function_242 neuron1577_1 (
      .a(input_layer[152]),
      .b(input_layer[909]),
      .c(~input_layer[573]),
      .d(input_layer[1300]),
      .e(input_layer[988]),
      .f(input_layer[1346]),
      .y(Y[1577]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1578_1
  function_167 neuron1578_1 (
      .a(input_layer[965]),
      .b(input_layer[203]),
      .c(input_layer[1247]),
      .d(~input_layer[983]),
      .e(input_layer[935]),
      .y(Y[1578]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_405 for neuron1579_1
  function_405 neuron1579_1 (
      .a(input_layer[196]),
      .b(~input_layer[1489]),
      .c(~input_layer[548]),
      .d(input_layer[891]),
      .e(~input_layer[1240]),
      .f(~input_layer[561]),
      .y(Y[1579]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1580_1
  function_120 neuron1580_1 (
      .a(input_layer[1308]),
      .b(~input_layer[694]),
      .c(input_layer[474]),
      .d(~input_layer[760]),
      .e(~input_layer[272]),
      .y(Y[1580]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1581_1
  function_4 neuron1581_1 (
      .a(input_layer[717]),
      .b(~input_layer[290]),
      .c(~input_layer[516]),
      .d(~input_layer[340]),
      .e(~input_layer[325]),
      .y(Y[1581]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1582_1
  function_11 neuron1582_1 (
      .a(~input_layer[1221]),
      .b(~input_layer[1250]),
      .c(input_layer[77]),
      .d(~input_layer[1338]),
      .y(Y[1582]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1583_1
  function_8 neuron1583_1 (
      .a(input_layer[251]),
      .b(input_layer[939]),
      .c(~input_layer[802]),
      .d(~input_layer[328]),
      .y(Y[1583]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1584_1
  function_47 neuron1584_1 (
      .a(input_layer[1417]),
      .b(input_layer[359]),
      .c(input_layer[1089]),
      .d(input_layer[84]),
      .e(input_layer[522]),
      .y(Y[1584]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1585_1
  function_95 neuron1585_1 (
      .a(input_layer[1165]),
      .b(~input_layer[584]),
      .c(~input_layer[83]),
      .d(~input_layer[669]),
      .y(Y[1585]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_377 for neuron1586_1
  function_377 neuron1586_1 (
      .a(~input_layer[720]),
      .b(~input_layer[772]),
      .c(input_layer[611]),
      .d(input_layer[1272]),
      .e(input_layer[895]),
      .f(input_layer[1452]),
      .y(Y[1586]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1587_1
  function_26 neuron1587_1 (
      .a(~input_layer[1164]),
      .y(Y[1587]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1588_1
  function_67 neuron1588_1 (
      .a(~input_layer[1001]),
      .b(~input_layer[1531]),
      .c(~input_layer[741]),
      .d(~input_layer[1160]),
      .e(~input_layer[1445]),
      .y(Y[1588]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1589_1
  function_12 neuron1589_1 (
      .a(input_layer[143]),
      .b(input_layer[771]),
      .c(~input_layer[1161]),
      .y(Y[1589]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1590_1
  function_89 neuron1590_1 (
      .a(input_layer[319]),
      .b(input_layer[812]),
      .c(~input_layer[455]),
      .d(~input_layer[1361]),
      .e(input_layer[1445]),
      .y(Y[1590]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1591_1
  function_8 neuron1591_1 (
      .a(input_layer[213]),
      .b(~input_layer[1264]),
      .c(input_layer[848]),
      .d(~input_layer[368]),
      .y(Y[1591]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1592_1
  function_12 neuron1592_1 (
      .a(input_layer[1476]),
      .b(~input_layer[415]),
      .c(~input_layer[1223]),
      .y(Y[1592]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1593_1
  function_16 neuron1593_1 (
      .a(input_layer[979]),
      .b(input_layer[760]),
      .y(Y[1593]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron1594_1
  function_183 neuron1594_1 (
      .a(~input_layer[1310]),
      .b(input_layer[631]),
      .c(input_layer[904]),
      .d(input_layer[369]),
      .e(input_layer[790]),
      .f(input_layer[232]),
      .y(Y[1594]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1595_1
  function_55 neuron1595_1 (
      .a(~input_layer[818]),
      .b(~input_layer[182]),
      .c(~input_layer[1382]),
      .d(~input_layer[1390]),
      .e(~input_layer[655]),
      .y(Y[1595]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron1596_1
  function_69 neuron1596_1 (
      .a(input_layer[817]),
      .b(~input_layer[542]),
      .c(~input_layer[439]),
      .d(input_layer[1323]),
      .e(input_layer[899]),
      .f(input_layer[1162]),
      .y(Y[1596]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1597_1
  function_97 neuron1597_1 (
      .a(~input_layer[467]),
      .b(~input_layer[322]),
      .c(~input_layer[1059]),
      .d(input_layer[182]),
      .e(~input_layer[788]),
      .y(Y[1597]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1598_1
  function_26 neuron1598_1 (
      .a(input_layer[800]),
      .y(Y[1598]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_200 for neuron1599_1
  function_200 neuron1599_1 (
      .a(~input_layer[775]),
      .b(input_layer[1052]),
      .c(input_layer[1245]),
      .d(~input_layer[650]),
      .e(~input_layer[809]),
      .f(input_layer[1250]),
      .y(Y[1599]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1600_1
  function_154 neuron1600_1 (
      .a(~input_layer[635]),
      .b(~input_layer[791]),
      .c(input_layer[1206]),
      .d(~input_layer[1001]),
      .e(input_layer[1255]),
      .f(input_layer[49]),
      .y(Y[1600]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1601_1
  function_0 neuron1601_1 (
      .a(~input_layer[1412]),
      .b(~input_layer[1319]),
      .c(input_layer[923]),
      .d(~input_layer[125]),
      .e(~input_layer[209]),
      .y(Y[1601]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1602_1
  function_100 neuron1602_1 (
      .a(~input_layer[412]),
      .b(input_layer[1425]),
      .c(~input_layer[1004]),
      .d(~input_layer[1330]),
      .e(input_layer[1469]),
      .f(~input_layer[774]),
      .y(Y[1602]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1603_1
  function_167 neuron1603_1 (
      .a(input_layer[1102]),
      .b(input_layer[1471]),
      .c(input_layer[1499]),
      .d(input_layer[300]),
      .e(~input_layer[619]),
      .y(Y[1603]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1604_1
  function_167 neuron1604_1 (
      .a(input_layer[661]),
      .b(~input_layer[591]),
      .c(input_layer[1114]),
      .d(input_layer[654]),
      .e(~input_layer[646]),
      .y(Y[1604]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1605_1
  function_42 neuron1605_1 (
      .a(input_layer[145]),
      .b(~input_layer[755]),
      .c(input_layer[1069]),
      .d(input_layer[241]),
      .y(Y[1605]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1606_1
  function_26 neuron1606_1 (
      .a(input_layer[1024]),
      .y(Y[1606]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1607_1
  function_26 neuron1607_1 (
      .a(input_layer[772]),
      .y(Y[1607]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_406 for neuron1608_1
  function_406 neuron1608_1 (
      .a(~input_layer[858]),
      .b(input_layer[571]),
      .c(~input_layer[1296]),
      .d(input_layer[836]),
      .e(input_layer[789]),
      .f(input_layer[592]),
      .y(Y[1608]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_389 for neuron1609_1
  function_389 neuron1609_1 (
      .a(input_layer[718]),
      .b(~input_layer[509]),
      .c(input_layer[1280]),
      .d(input_layer[1266]),
      .e(input_layer[158]),
      .f(input_layer[284]),
      .y(Y[1609]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron1610_1
  function_75 neuron1610_1 (
      .a(~input_layer[688]),
      .b(~input_layer[635]),
      .c(input_layer[677]),
      .d(input_layer[1296]),
      .e(input_layer[458]),
      .y(Y[1610]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_407 for neuron1611_1
  function_407 neuron1611_1 (
      .a(~input_layer[1320]),
      .b(~input_layer[1186]),
      .c(input_layer[1293]),
      .d(~input_layer[430]),
      .e(input_layer[1228]),
      .f(input_layer[766]),
      .y(Y[1611]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1612_1
  function_35 neuron1612_1 (
      .a(~input_layer[1369]),
      .b(~input_layer[457]),
      .c(~input_layer[1529]),
      .d(input_layer[599]),
      .e(input_layer[1090]),
      .y(Y[1612]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1613_1
  function_271 neuron1613_1 (
      .a(input_layer[813]),
      .b(~input_layer[1191]),
      .c(input_layer[1548]),
      .d(input_layer[680]),
      .e(input_layer[219]),
      .y(Y[1613]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1614_1
  function_8 neuron1614_1 (
      .a(input_layer[634]),
      .b(input_layer[550]),
      .c(~input_layer[1170]),
      .d(input_layer[716]),
      .y(Y[1614]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1615_1
  function_47 neuron1615_1 (
      .a(input_layer[972]),
      .b(input_layer[238]),
      .c(input_layer[151]),
      .d(input_layer[1414]),
      .e(input_layer[1060]),
      .y(Y[1615]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1616_1
  function_27 neuron1616_1 (
      .a(input_layer[325]),
      .b(~input_layer[459]),
      .c(~input_layer[861]),
      .y(Y[1616]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1617_1
  function_26 neuron1617_1 (
      .a(input_layer[913]),
      .y(Y[1617]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1618_1
  function_8 neuron1618_1 (
      .a(input_layer[1332]),
      .b(input_layer[662]),
      .c(input_layer[1107]),
      .d(~input_layer[465]),
      .y(Y[1618]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_408 for neuron1619_1
  function_408 neuron1619_1 (
      .a(input_layer[1475]),
      .b(~input_layer[1242]),
      .c(input_layer[739]),
      .d(input_layer[1424]),
      .e(input_layer[659]),
      .f(input_layer[706]),
      .y(Y[1619]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1620_1
  function_334 neuron1620_1 (
      .a(~input_layer[1218]),
      .b(~input_layer[350]),
      .c(input_layer[655]),
      .d(input_layer[72]),
      .e(input_layer[98]),
      .y(Y[1620]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1621_1
  function_97 neuron1621_1 (
      .a(~input_layer[1049]),
      .b(input_layer[923]),
      .c(~input_layer[1002]),
      .d(~input_layer[973]),
      .e(~input_layer[324]),
      .y(Y[1621]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1622_1
  function_8 neuron1622_1 (
      .a(input_layer[1002]),
      .b(~input_layer[934]),
      .c(input_layer[849]),
      .d(~input_layer[1104]),
      .y(Y[1622]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1623_1
  function_29 neuron1623_1 (
      .a(~input_layer[981]),
      .b(input_layer[1255]),
      .y(Y[1623]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1624_1
  function_128 neuron1624_1 (
      .a(input_layer[1254]),
      .b(~input_layer[802]),
      .c(input_layer[1269]),
      .d(input_layer[808]),
      .y(Y[1624]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1625_1
  function_1 neuron1625_1 (
      .a(~input_layer[805]),
      .b(input_layer[681]),
      .c(~input_layer[1270]),
      .d(~input_layer[268]),
      .y(Y[1625]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1626_1
  function_67 neuron1626_1 (
      .a(~input_layer[195]),
      .b(~input_layer[832]),
      .c(~input_layer[436]),
      .d(~input_layer[508]),
      .e(~input_layer[562]),
      .y(Y[1626]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1627_1
  function_17 neuron1627_1 (
      .a(input_layer[1221]),
      .b(input_layer[1545]),
      .c(~input_layer[1304]),
      .y(Y[1627]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1628_1
  function_298 neuron1628_1 (
      .a(~input_layer[754]),
      .b(~input_layer[1241]),
      .c(~input_layer[241]),
      .d(input_layer[667]),
      .e(~input_layer[519]),
      .f(input_layer[534]),
      .y(Y[1628]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_409 for neuron1629_1
  function_409 neuron1629_1 (
      .a(~input_layer[1170]),
      .b(~input_layer[778]),
      .c(input_layer[1181]),
      .d(~input_layer[769]),
      .e(input_layer[1193]),
      .f(~input_layer[870]),
      .y(Y[1629]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1630_1
  function_42 neuron1630_1 (
      .a(input_layer[290]),
      .b(input_layer[904]),
      .c(input_layer[1336]),
      .d(input_layer[87]),
      .y(Y[1630]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_285 for neuron1631_1
  function_285 neuron1631_1 (
      .a(~input_layer[1057]),
      .b(~input_layer[970]),
      .c(~input_layer[265]),
      .d(input_layer[788]),
      .e(input_layer[421]),
      .f(input_layer[340]),
      .y(Y[1631]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1632_1
  function_107 neuron1632_1 (
      .a(~input_layer[1362]),
      .b(~input_layer[82]),
      .c(~input_layer[1555]),
      .d(input_layer[617]),
      .e(input_layer[1267]),
      .y(Y[1632]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1633_1
  function_87 neuron1633_1 (
      .a(input_layer[924]),
      .b(~input_layer[591]),
      .c(input_layer[73]),
      .d(~input_layer[844]),
      .e(input_layer[609]),
      .y(Y[1633]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_410 for neuron1634_1
  function_410 neuron1634_1 (
      .a(~input_layer[911]),
      .b(~input_layer[244]),
      .c(~input_layer[1191]),
      .d(input_layer[934]),
      .e(~input_layer[241]),
      .f(input_layer[653]),
      .y(Y[1634]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1635_1
  function_49 neuron1635_1 (
      .a(~input_layer[382]),
      .b(input_layer[825]),
      .c(~input_layer[515]),
      .d(~input_layer[648]),
      .e(input_layer[1469]),
      .y(Y[1635]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1636_1
  function_39 neuron1636_1 (
      .a(~input_layer[261]),
      .b(input_layer[438]),
      .c(~input_layer[1040]),
      .y(Y[1636]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron1637_1
  function_145 neuron1637_1 (
      .a(input_layer[1280]),
      .b(~input_layer[1072]),
      .c(~input_layer[877]),
      .d(input_layer[94]),
      .e(input_layer[271]),
      .y(Y[1637]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_411 for neuron1638_1
  function_411 neuron1638_1 (
      .a(~input_layer[530]),
      .b(input_layer[1543]),
      .c(input_layer[486]),
      .d(input_layer[81]),
      .e(~input_layer[1262]),
      .f(input_layer[1179]),
      .y(Y[1638]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1639_1
  function_3 neuron1639_1 (
      .a(~input_layer[187]),
      .b(~input_layer[697]),
      .c(~input_layer[644]),
      .d(~input_layer[668]),
      .y(Y[1639]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_300 for neuron1640_1
  function_300 neuron1640_1 (
      .a(input_layer[1421]),
      .b(~input_layer[206]),
      .c(~input_layer[1255]),
      .d(input_layer[1057]),
      .e(input_layer[518]),
      .y(Y[1640]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1641_1
  function_97 neuron1641_1 (
      .a(input_layer[385]),
      .b(~input_layer[84]),
      .c(~input_layer[458]),
      .d(~input_layer[1408]),
      .e(~input_layer[1055]),
      .y(Y[1641]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1642_1
  function_4 neuron1642_1 (
      .a(input_layer[1266]),
      .b(~input_layer[1353]),
      .c(~input_layer[674]),
      .d(~input_layer[781]),
      .e(~input_layer[163]),
      .y(Y[1642]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1643_1
  function_48 neuron1643_1 (
      .a(input_layer[354]),
      .b(input_layer[941]),
      .c(input_layer[947]),
      .d(input_layer[1220]),
      .e(~input_layer[1430]),
      .y(Y[1643]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_412 for neuron1644_1
  function_412 neuron1644_1 (
      .a(~input_layer[628]),
      .b(input_layer[1241]),
      .c(~input_layer[528]),
      .d(input_layer[893]),
      .e(~input_layer[981]),
      .y(Y[1644]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1645_1
  function_24 neuron1645_1 (
      .a(~input_layer[1056]),
      .b(~input_layer[247]),
      .c(input_layer[325]),
      .y(Y[1645]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1646_1
  function_16 neuron1646_1 (
      .a(input_layer[557]),
      .b(~input_layer[1388]),
      .y(Y[1646]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1647_1
  function_87 neuron1647_1 (
      .a(input_layer[255]),
      .b(~input_layer[1540]),
      .c(input_layer[848]),
      .d(input_layer[694]),
      .e(~input_layer[983]),
      .y(Y[1647]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1648_1
  function_27 neuron1648_1 (
      .a(~input_layer[442]),
      .b(input_layer[647]),
      .c(~input_layer[1535]),
      .y(Y[1648]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1649_1
  function_67 neuron1649_1 (
      .a(~input_layer[513]),
      .b(~input_layer[739]),
      .c(~input_layer[1222]),
      .d(~input_layer[180]),
      .e(input_layer[1305]),
      .y(Y[1649]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_413 for neuron1650_1
  function_413 neuron1650_1 (
      .a(~input_layer[977]),
      .b(~input_layer[148]),
      .c(input_layer[1353]),
      .d(input_layer[1360]),
      .e(input_layer[1369]),
      .f(input_layer[549]),
      .y(Y[1650]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_414 for neuron1651_1
  function_414 neuron1651_1 (
      .a(~input_layer[825]),
      .b(~input_layer[800]),
      .c(input_layer[598]),
      .d(~input_layer[1354]),
      .e(~input_layer[224]),
      .f(~input_layer[1452]),
      .y(Y[1651]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1652] = 1'b0;

  // instantiate function_415 for neuron1653_1
  function_415 neuron1653_1 (
      .a(~input_layer[748]),
      .b(~input_layer[611]),
      .c(input_layer[1051]),
      .d(~input_layer[1501]),
      .e(input_layer[865]),
      .f(input_layer[1154]),
      .y(Y[1653]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1654_1
  function_16 neuron1654_1 (
      .a(~input_layer[366]),
      .b(input_layer[1061]),
      .y(Y[1654]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1655_1
  function_154 neuron1655_1 (
      .a(~input_layer[138]),
      .b(~input_layer[751]),
      .c(~input_layer[853]),
      .d(input_layer[1413]),
      .e(~input_layer[284]),
      .f(~input_layer[1178]),
      .y(Y[1655]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1656_1
  function_16 neuron1656_1 (
      .a(input_layer[1029]),
      .b(input_layer[830]),
      .y(Y[1656]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1657_1
  function_214 neuron1657_1 (
      .a(input_layer[328]),
      .b(input_layer[152]),
      .c(input_layer[566]),
      .d(input_layer[490]),
      .e(~input_layer[534]),
      .f(~input_layer[627]),
      .y(Y[1657]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_416 for neuron1658_1
  function_416 neuron1658_1 (
      .a(input_layer[1247]),
      .b(input_layer[455]),
      .c(~input_layer[1142]),
      .d(~input_layer[82]),
      .e(~input_layer[262]),
      .f(~input_layer[988]),
      .y(Y[1658]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron1659_1
  function_221 neuron1659_1 (
      .a(input_layer[1170]),
      .b(input_layer[322]),
      .c(~input_layer[297]),
      .d(~input_layer[289]),
      .e(input_layer[765]),
      .f(input_layer[163]),
      .y(Y[1659]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_320 for neuron1660_1
  function_320 neuron1660_1 (
      .a(input_layer[808]),
      .b(input_layer[1390]),
      .c(~input_layer[598]),
      .d(input_layer[1337]),
      .e(~input_layer[1202]),
      .f(input_layer[431]),
      .y(Y[1660]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1661] = 1'b0;

  // instantiate function_241 for neuron1662_1
  function_241 neuron1662_1 (
      .a(input_layer[1059]),
      .b(input_layer[942]),
      .c(input_layer[82]),
      .d(~input_layer[399]),
      .e(~input_layer[1376]),
      .f(input_layer[899]),
      .y(Y[1662]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1663_1
  function_47 neuron1663_1 (
      .a(input_layer[1469]),
      .b(input_layer[737]),
      .c(input_layer[1555]),
      .d(input_layer[1524]),
      .e(~input_layer[643]),
      .y(Y[1663]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_396 for neuron1664_1
  function_396 neuron1664_1 (
      .a(input_layer[190]),
      .b(input_layer[86]),
      .c(~input_layer[1038]),
      .d(~input_layer[351]),
      .e(~input_layer[232]),
      .y(Y[1664]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1665_1
  function_29 neuron1665_1 (
      .a(~input_layer[1043]),
      .b(~input_layer[1335]),
      .y(Y[1665]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_417 for neuron1666_1
  function_417 neuron1666_1 (
      .a(~input_layer[652]),
      .b(~input_layer[709]),
      .c(~input_layer[202]),
      .d(input_layer[583]),
      .e(~input_layer[1084]),
      .f(input_layer[1156]),
      .y(Y[1666]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1667_1
  function_30 neuron1667_1 (
      .a(input_layer[790]),
      .b(input_layer[1087]),
      .c(~input_layer[998]),
      .d(~input_layer[1186]),
      .y(Y[1667]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron1668_1
  function_13 neuron1668_1 (
      .a(~input_layer[1102]),
      .b(input_layer[623]),
      .c(~input_layer[1057]),
      .d(~input_layer[93]),
      .y(Y[1668]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1669_1
  function_12 neuron1669_1 (
      .a(input_layer[860]),
      .b(~input_layer[1147]),
      .c(~input_layer[266]),
      .y(Y[1669]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_418 for neuron1670_1
  function_418 neuron1670_1 (
      .a(input_layer[709]),
      .b(~input_layer[308]),
      .c(~input_layer[1020]),
      .d(~input_layer[1000]),
      .e(~input_layer[1198]),
      .y(Y[1670]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1671_1
  function_24 neuron1671_1 (
      .a(input_layer[385]),
      .b(~input_layer[999]),
      .c(~input_layer[1390]),
      .y(Y[1671]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_369 for neuron1672_1
  function_369 neuron1672_1 (
      .a(~input_layer[536]),
      .b(input_layer[771]),
      .c(~input_layer[1004]),
      .d(~input_layer[949]),
      .e(input_layer[249]),
      .f(input_layer[945]),
      .y(Y[1672]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1673_1
  function_60 neuron1673_1 (
      .a(input_layer[464]),
      .b(input_layer[1429]),
      .c(input_layer[304]),
      .d(input_layer[485]),
      .e(input_layer[64]),
      .y(Y[1673]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1674_1
  function_28 neuron1674_1 (
      .a(~input_layer[496]),
      .b(~input_layer[886]),
      .c(~input_layer[1001]),
      .d(~input_layer[1295]),
      .e(~input_layer[1226]),
      .f(~input_layer[604]),
      .y(Y[1674]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_313 for neuron1675_1
  function_313 neuron1675_1 (
      .a(~input_layer[495]),
      .b(input_layer[1408]),
      .c(~input_layer[1265]),
      .d(~input_layer[751]),
      .e(input_layer[338]),
      .f(input_layer[729]),
      .y(Y[1675]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1676_1
  function_107 neuron1676_1 (
      .a(~input_layer[422]),
      .b(~input_layer[1244]),
      .c(~input_layer[1048]),
      .d(input_layer[338]),
      .e(input_layer[1505]),
      .y(Y[1676]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_136 for neuron1677_1
  function_136 neuron1677_1 (
      .a(input_layer[1370]),
      .b(~input_layer[187]),
      .c(input_layer[1309]),
      .d(input_layer[269]),
      .e(input_layer[1560]),
      .f(input_layer[127]),
      .y(Y[1677]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1678_1
  function_16 neuron1678_1 (
      .a(input_layer[610]),
      .b(input_layer[589]),
      .y(Y[1678]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1679_1
  function_46 neuron1679_1 (
      .a(input_layer[698]),
      .b(input_layer[777]),
      .c(~input_layer[1194]),
      .d(input_layer[888]),
      .e(input_layer[376]),
      .y(Y[1679]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_419 for neuron1680_1
  function_419 neuron1680_1 (
      .a(input_layer[1542]),
      .b(~input_layer[880]),
      .c(~input_layer[273]),
      .d(~input_layer[910]),
      .e(~input_layer[88]),
      .f(input_layer[1067]),
      .y(Y[1680]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_420 for neuron1681_1
  function_420 neuron1681_1 (
      .a(input_layer[642]),
      .b(~input_layer[245]),
      .c(~input_layer[412]),
      .d(input_layer[757]),
      .e(input_layer[898]),
      .f(~input_layer[1197]),
      .y(Y[1681]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1682_1
  function_149 neuron1682_1 (
      .a(~input_layer[265]),
      .b(input_layer[716]),
      .c(~input_layer[593]),
      .d(input_layer[610]),
      .y(Y[1682]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_329 for neuron1683_1
  function_329 neuron1683_1 (
      .a(input_layer[529]),
      .b(~input_layer[853]),
      .c(~input_layer[74]),
      .d(~input_layer[416]),
      .e(input_layer[1146]),
      .f(input_layer[785]),
      .y(Y[1683]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1684_1
  function_48 neuron1684_1 (
      .a(input_layer[973]),
      .b(input_layer[139]),
      .c(input_layer[861]),
      .d(input_layer[80]),
      .e(input_layer[1244]),
      .y(Y[1684]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_421 for neuron1685_1
  function_421 neuron1685_1 (
      .a(~input_layer[435]),
      .b(input_layer[134]),
      .c(~input_layer[961]),
      .d(~input_layer[991]),
      .e(input_layer[1149]),
      .f(input_layer[865]),
      .y(Y[1685]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron1686_1
  function_82 neuron1686_1 (
      .a(~input_layer[775]),
      .b(~input_layer[662]),
      .c(~input_layer[86]),
      .d(input_layer[520]),
      .e(input_layer[1110]),
      .f(~input_layer[56]),
      .y(Y[1686]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron1687_1
  function_36 neuron1687_1 (
      .a(input_layer[1219]),
      .b(input_layer[605]),
      .c(input_layer[1155]),
      .d(input_layer[1277]),
      .e(input_layer[360]),
      .f(input_layer[1306]),
      .y(Y[1687]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_349 for neuron1688_1
  function_349 neuron1688_1 (
      .a(input_layer[595]),
      .b(input_layer[622]),
      .c(~input_layer[971]),
      .d(~input_layer[156]),
      .e(input_layer[796]),
      .y(Y[1688]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_71 for neuron1689_1
  function_71 neuron1689_1 (
      .a(input_layer[1486]),
      .b(input_layer[142]),
      .c(~input_layer[1246]),
      .d(~input_layer[416]),
      .e(input_layer[959]),
      .f(input_layer[236]),
      .y(Y[1689]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1690_1
  function_67 neuron1690_1 (
      .a(~input_layer[881]),
      .b(~input_layer[746]),
      .c(~input_layer[849]),
      .d(~input_layer[1245]),
      .e(~input_layer[540]),
      .y(Y[1690]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1691_1
  function_3 neuron1691_1 (
      .a(~input_layer[1056]),
      .b(~input_layer[1109]),
      .c(~input_layer[298]),
      .d(~input_layer[1161]),
      .y(Y[1691]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1692_1
  function_128 neuron1692_1 (
      .a(~input_layer[529]),
      .b(~input_layer[721]),
      .c(~input_layer[377]),
      .d(input_layer[955]),
      .y(Y[1692]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1693_1
  function_12 neuron1693_1 (
      .a(input_layer[1379]),
      .b(~input_layer[213]),
      .c(input_layer[588]),
      .y(Y[1693]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1694] = 1'b1;

  // instantiate function_8 for neuron1695_1
  function_8 neuron1695_1 (
      .a(input_layer[941]),
      .b(input_layer[1421]),
      .c(input_layer[827]),
      .d(input_layer[989]),
      .y(Y[1695]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1696_1
  function_24 neuron1696_1 (
      .a(~input_layer[585]),
      .b(~input_layer[775]),
      .c(input_layer[178]),
      .y(Y[1696]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1697_1
  function_48 neuron1697_1 (
      .a(input_layer[198]),
      .b(input_layer[927]),
      .c(~input_layer[319]),
      .d(input_layer[79]),
      .e(~input_layer[1139]),
      .y(Y[1697]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1698_1
  function_106 neuron1698_1 (
      .a(input_layer[1247]),
      .b(~input_layer[1417]),
      .c(~input_layer[1320]),
      .d(input_layer[1294]),
      .y(Y[1698]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1699_1
  function_29 neuron1699_1 (
      .a(~input_layer[713]),
      .b(~input_layer[906]),
      .y(Y[1699]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1700_1
  function_29 neuron1700_1 (
      .a(~input_layer[989]),
      .b(~input_layer[488]),
      .y(Y[1700]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1701_1
  function_27 neuron1701_1 (
      .a(~input_layer[908]),
      .b(~input_layer[873]),
      .c(~input_layer[1417]),
      .y(Y[1701]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_420 for neuron1702_1
  function_420 neuron1702_1 (
      .a(~input_layer[1246]),
      .b(~input_layer[1015]),
      .c(input_layer[1096]),
      .d(input_layer[148]),
      .e(~input_layer[795]),
      .f(input_layer[889]),
      .y(Y[1702]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1703_1
  function_29 neuron1703_1 (
      .a(~input_layer[755]),
      .b(~input_layer[153]),
      .y(Y[1703]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_422 for neuron1704_1
  function_422 neuron1704_1 (
      .a(input_layer[497]),
      .b(input_layer[1056]),
      .c(input_layer[1144]),
      .d(~input_layer[1254]),
      .e(~input_layer[1415]),
      .f(~input_layer[452]),
      .y(Y[1704]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1705_1
  function_113 neuron1705_1 (
      .a(~input_layer[702]),
      .b(~input_layer[696]),
      .c(input_layer[82]),
      .d(input_layer[997]),
      .e(~input_layer[1356]),
      .y(Y[1705]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1706_1
  function_31 neuron1706_1 (
      .a(~input_layer[870]),
      .b(~input_layer[820]),
      .c(input_layer[882]),
      .d(input_layer[1148]),
      .y(Y[1706]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1707_1
  function_29 neuron1707_1 (
      .a(~input_layer[1087]),
      .b(~input_layer[1080]),
      .y(Y[1707]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1708_1
  function_186 neuron1708_1 (
      .a(input_layer[1493]),
      .b(input_layer[1353]),
      .c(~input_layer[192]),
      .d(~input_layer[126]),
      .y(Y[1708]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1709_1
  function_78 neuron1709_1 (
      .a(~input_layer[302]),
      .b(~input_layer[962]),
      .c(~input_layer[999]),
      .d(~input_layer[964]),
      .e(~input_layer[1338]),
      .f(input_layer[121]),
      .y(Y[1709]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron1710_1
  function_121 neuron1710_1 (
      .a(input_layer[1435]),
      .b(~input_layer[998]),
      .c(input_layer[95]),
      .d(input_layer[1551]),
      .e(input_layer[390]),
      .y(Y[1710]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1711_1
  function_123 neuron1711_1 (
      .a(input_layer[812]),
      .b(input_layer[188]),
      .c(input_layer[1085]),
      .d(~input_layer[1039]),
      .y(Y[1711]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1712_1
  function_17 neuron1712_1 (
      .a(input_layer[1480]),
      .b(input_layer[1140]),
      .c(input_layer[1423]),
      .y(Y[1712]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1713_1
  function_123 neuron1713_1 (
      .a(input_layer[1070]),
      .b(input_layer[478]),
      .c(~input_layer[1274]),
      .d(~input_layer[851]),
      .y(Y[1713]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1714] = 1'b0;

  // instantiate function_155 for neuron1715_1
  function_155 neuron1715_1 (
      .a(~input_layer[134]),
      .b(~input_layer[835]),
      .c(~input_layer[1354]),
      .d(input_layer[1390]),
      .e(input_layer[1448]),
      .f(~input_layer[1063]),
      .y(Y[1715]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1716_1
  function_271 neuron1716_1 (
      .a(input_layer[1127]),
      .b(input_layer[789]),
      .c(~input_layer[1198]),
      .d(~input_layer[750]),
      .e(~input_layer[332]),
      .y(Y[1716]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_423 for neuron1717_1
  function_423 neuron1717_1 (
      .a(input_layer[861]),
      .b(~input_layer[1035]),
      .c(input_layer[1192]),
      .d(~input_layer[1280]),
      .e(input_layer[666]),
      .f(~input_layer[1551]),
      .y(Y[1717]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1718_1
  function_113 neuron1718_1 (
      .a(~input_layer[918]),
      .b(input_layer[1293]),
      .c(~input_layer[945]),
      .d(~input_layer[1025]),
      .e(input_layer[451]),
      .y(Y[1718]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1719_1
  function_0 neuron1719_1 (
      .a(~input_layer[136]),
      .b(~input_layer[1137]),
      .c(~input_layer[1540]),
      .d(input_layer[979]),
      .e(~input_layer[216]),
      .y(Y[1719]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1720_1
  function_67 neuron1720_1 (
      .a(~input_layer[909]),
      .b(~input_layer[516]),
      .c(~input_layer[249]),
      .d(~input_layer[893]),
      .e(~input_layer[511]),
      .y(Y[1720]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_424 for neuron1721_1
  function_424 neuron1721_1 (
      .a(input_layer[919]),
      .b(~input_layer[1246]),
      .c(~input_layer[345]),
      .d(input_layer[965]),
      .e(input_layer[1004]),
      .f(~input_layer[446]),
      .y(Y[1721]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1722_1
  function_87 neuron1722_1 (
      .a(input_layer[510]),
      .b(~input_layer[1125]),
      .c(input_layer[1558]),
      .d(input_layer[104]),
      .e(input_layer[4]),
      .y(Y[1722]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1723_1
  function_27 neuron1723_1 (
      .a(~input_layer[1482]),
      .b(~input_layer[1354]),
      .c(input_layer[79]),
      .y(Y[1723]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1724_1
  function_149 neuron1724_1 (
      .a(~input_layer[1364]),
      .b(~input_layer[1257]),
      .c(input_layer[1237]),
      .d(~input_layer[137]),
      .y(Y[1724]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1725_1
  function_92 neuron1725_1 (
      .a(input_layer[1057]),
      .b(input_layer[1019]),
      .c(input_layer[890]),
      .d(input_layer[1142]),
      .e(input_layer[1106]),
      .f(~input_layer[1406]),
      .y(Y[1725]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron1726_1
  function_84 neuron1726_1 (
      .a(~input_layer[913]),
      .b(input_layer[352]),
      .c(input_layer[312]),
      .d(input_layer[1204]),
      .e(~input_layer[1502]),
      .y(Y[1726]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1727_1
  function_26 neuron1727_1 (
      .a(input_layer[196]),
      .y(Y[1727]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_233 for neuron1728_1
  function_233 neuron1728_1 (
      .a(input_layer[816]),
      .b(input_layer[1383]),
      .c(~input_layer[232]),
      .d(~input_layer[431]),
      .e(~input_layer[64]),
      .f(input_layer[1399]),
      .y(Y[1728]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_425 for neuron1729_1
  function_425 neuron1729_1 (
      .a(input_layer[631]),
      .b(input_layer[1541]),
      .c(input_layer[1323]),
      .d(~input_layer[1192]),
      .e(~input_layer[1193]),
      .f(~input_layer[404]),
      .y(Y[1729]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1730_1
  function_35 neuron1730_1 (
      .a(~input_layer[1143]),
      .b(~input_layer[1101]),
      .c(~input_layer[148]),
      .d(~input_layer[431]),
      .e(~input_layer[358]),
      .y(Y[1730]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1731_1
  function_87 neuron1731_1 (
      .a(input_layer[463]),
      .b(~input_layer[1255]),
      .c(input_layer[821]),
      .d(input_layer[1525]),
      .e(~input_layer[995]),
      .y(Y[1731]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron1732_1
  function_62 neuron1732_1 (
      .a(input_layer[621]),
      .b(~input_layer[761]),
      .c(input_layer[993]),
      .d(input_layer[1069]),
      .e(input_layer[677]),
      .f(~input_layer[657]),
      .y(Y[1732]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_23 for neuron1733_1
  function_23 neuron1733_1 (
      .a(input_layer[1170]),
      .b(~input_layer[1156]),
      .c(~input_layer[1306]),
      .d(~input_layer[1542]),
      .e(~input_layer[27]),
      .f(~input_layer[24]),
      .y(Y[1733]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron1734_1
  function_210 neuron1734_1 (
      .a(~input_layer[1480]),
      .b(input_layer[911]),
      .c(~input_layer[621]),
      .d(~input_layer[837]),
      .e(~input_layer[1533]),
      .f(input_layer[597]),
      .y(Y[1734]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1735_1
  function_99 neuron1735_1 (
      .a(input_layer[1135]),
      .b(input_layer[442]),
      .c(input_layer[379]),
      .d(~input_layer[860]),
      .e(~input_layer[80]),
      .y(Y[1735]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1736_1
  function_27 neuron1736_1 (
      .a(~input_layer[776]),
      .b(~input_layer[551]),
      .c(input_layer[425]),
      .y(Y[1736]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1737_1
  function_56 neuron1737_1 (
      .a(~input_layer[976]),
      .b(input_layer[271]),
      .c(~input_layer[193]),
      .d(input_layer[844]),
      .e(~input_layer[26]),
      .y(Y[1737]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1738_1
  function_46 neuron1738_1 (
      .a(input_layer[1199]),
      .b(input_layer[569]),
      .c(input_layer[233]),
      .d(input_layer[1123]),
      .e(input_layer[1032]),
      .y(Y[1738]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1739_1
  function_17 neuron1739_1 (
      .a(input_layer[754]),
      .b(input_layer[906]),
      .c(input_layer[79]),
      .y(Y[1739]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_198 for neuron1740_1
  function_198 neuron1740_1 (
      .a(input_layer[1312]),
      .b(~input_layer[210]),
      .c(~input_layer[912]),
      .d(~input_layer[1447]),
      .e(input_layer[359]),
      .f(input_layer[311]),
      .y(Y[1740]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_86 for neuron1741_1
  function_86 neuron1741_1 (
      .a(input_layer[1077]),
      .b(input_layer[241]),
      .c(input_layer[200]),
      .d(input_layer[974]),
      .e(input_layer[1426]),
      .f(~input_layer[99]),
      .y(Y[1741]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1742_1
  function_167 neuron1742_1 (
      .a(input_layer[197]),
      .b(input_layer[611]),
      .c(input_layer[438]),
      .d(~input_layer[1547]),
      .e(input_layer[909]),
      .y(Y[1742]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1743_1
  function_92 neuron1743_1 (
      .a(input_layer[304]),
      .b(~input_layer[319]),
      .c(input_layer[307]),
      .d(~input_layer[474]),
      .e(~input_layer[368]),
      .f(~input_layer[55]),
      .y(Y[1743]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_426 for neuron1744_1
  function_426 neuron1744_1 (
      .a(input_layer[490]),
      .b(~input_layer[565]),
      .c(~input_layer[1430]),
      .d(~input_layer[457]),
      .e(input_layer[232]),
      .f(input_layer[1561]),
      .y(Y[1744]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1745_1
  function_19 neuron1745_1 (
      .a(~input_layer[1075]),
      .b(~input_layer[1236]),
      .c(input_layer[987]),
      .d(input_layer[516]),
      .y(Y[1745]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_212 for neuron1746_1
  function_212 neuron1746_1 (
      .a(~input_layer[1323]),
      .b(input_layer[485]),
      .c(input_layer[215]),
      .d(input_layer[1271]),
      .e(~input_layer[1303]),
      .y(Y[1746]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_275 for neuron1747_1
  function_275 neuron1747_1 (
      .a(input_layer[138]),
      .b(~input_layer[942]),
      .c(input_layer[790]),
      .d(input_layer[1365]),
      .e(input_layer[932]),
      .f(input_layer[505]),
      .y(Y[1747]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1748_1
  function_7 neuron1748_1 (
      .a(input_layer[543]),
      .b(~input_layer[207]),
      .c(input_layer[1469]),
      .d(~input_layer[252]),
      .y(Y[1748]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_257 for neuron1749_1
  function_257 neuron1749_1 (
      .a(input_layer[553]),
      .b(input_layer[1332]),
      .c(input_layer[1387]),
      .d(~input_layer[936]),
      .e(~input_layer[349]),
      .f(~input_layer[288]),
      .y(Y[1749]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1750_1
  function_11 neuron1750_1 (
      .a(~input_layer[1271]),
      .b(input_layer[541]),
      .c(input_layer[95]),
      .d(~input_layer[1284]),
      .y(Y[1750]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1751_1
  function_26 neuron1751_1 (
      .a(~input_layer[205]),
      .y(Y[1751]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1752_1
  function_100 neuron1752_1 (
      .a(~input_layer[1419]),
      .b(~input_layer[181]),
      .c(~input_layer[335]),
      .d(input_layer[1394]),
      .e(~input_layer[284]),
      .f(~input_layer[42]),
      .y(Y[1752]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_427 for neuron1753_1
  function_427 neuron1753_1 (
      .a(input_layer[1138]),
      .b(~input_layer[1422]),
      .c(~input_layer[511]),
      .d(~input_layer[566]),
      .e(input_layer[402]),
      .f(~input_layer[102]),
      .y(Y[1753]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_428 for neuron1754_1
  function_428 neuron1754_1 (
      .a(input_layer[970]),
      .b(input_layer[152]),
      .c(~input_layer[409]),
      .d(~input_layer[1042]),
      .e(~input_layer[360]),
      .f(input_layer[1330]),
      .y(Y[1754]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1755_1
  function_16 neuron1755_1 (
      .a(input_layer[353]),
      .b(input_layer[243]),
      .y(Y[1755]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1756_1
  function_330 neuron1756_1 (
      .a(~input_layer[365]),
      .b(input_layer[776]),
      .c(~input_layer[316]),
      .d(~input_layer[1139]),
      .e(~input_layer[834]),
      .y(Y[1756]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1757_1
  function_44 neuron1757_1 (
      .a(~input_layer[246]),
      .b(~input_layer[515]),
      .c(input_layer[1529]),
      .d(input_layer[1436]),
      .e(input_layer[1095]),
      .y(Y[1757]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1758_1
  function_29 neuron1758_1 (
      .a(~input_layer[711]),
      .b(~input_layer[572]),
      .y(Y[1758]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1759_1
  function_67 neuron1759_1 (
      .a(~input_layer[940]),
      .b(input_layer[1190]),
      .c(~input_layer[1470]),
      .d(~input_layer[1355]),
      .e(~input_layer[96]),
      .y(Y[1759]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1760_1
  function_29 neuron1760_1 (
      .a(~input_layer[687]),
      .b(input_layer[411]),
      .y(Y[1760]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1761_1
  function_120 neuron1761_1 (
      .a(input_layer[808]),
      .b(input_layer[1031]),
      .c(~input_layer[1475]),
      .d(~input_layer[873]),
      .e(input_layer[230]),
      .y(Y[1761]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1762_1
  function_0 neuron1762_1 (
      .a(~input_layer[694]),
      .b(~input_layer[1433]),
      .c(~input_layer[573]),
      .d(input_layer[980]),
      .e(~input_layer[249]),
      .y(Y[1762]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1763_1
  function_26 neuron1763_1 (
      .a(input_layer[1147]),
      .y(Y[1763]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1764_1
  function_76 neuron1764_1 (
      .a(input_layer[816]),
      .b(input_layer[149]),
      .c(input_layer[949]),
      .d(input_layer[237]),
      .e(input_layer[506]),
      .f(~input_layer[427]),
      .y(Y[1764]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron1765_1
  function_70 neuron1765_1 (
      .a(~input_layer[200]),
      .b(input_layer[433]),
      .c(~input_layer[1337]),
      .d(~input_layer[1329]),
      .e(~input_layer[1500]),
      .f(~input_layer[101]),
      .y(Y[1765]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1766_1
  function_29 neuron1766_1 (
      .a(~input_layer[1478]),
      .b(input_layer[466]),
      .y(Y[1766]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1767_1
  function_27 neuron1767_1 (
      .a(input_layer[602]),
      .b(input_layer[1314]),
      .c(~input_layer[1168]),
      .y(Y[1767]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_338 for neuron1768_1
  function_338 neuron1768_1 (
      .a(input_layer[264]),
      .b(input_layer[1331]),
      .c(~input_layer[1378]),
      .d(input_layer[871]),
      .e(~input_layer[1473]),
      .f(~input_layer[468]),
      .y(Y[1768]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1769_1
  function_17 neuron1769_1 (
      .a(input_layer[1241]),
      .b(input_layer[564]),
      .c(input_layer[310]),
      .y(Y[1769]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1770_1
  function_29 neuron1770_1 (
      .a(~input_layer[475]),
      .b(~input_layer[1026]),
      .y(Y[1770]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron1771_1
  function_74 neuron1771_1 (
      .a(~input_layer[1494]),
      .b(~input_layer[1095]),
      .c(input_layer[766]),
      .d(~input_layer[88]),
      .e(input_layer[1]),
      .f(input_layer[115]),
      .y(Y[1771]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_22 for neuron1772_1
  function_22 neuron1772_1 (
      .a(input_layer[1018]),
      .b(~input_layer[977]),
      .c(~input_layer[811]),
      .d(input_layer[1207]),
      .e(input_layer[1363]),
      .f(~input_layer[122]),
      .y(Y[1772]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_429 for neuron1773_1
  function_429 neuron1773_1 (
      .a(~input_layer[981]),
      .b(~input_layer[76]),
      .c(input_layer[1329]),
      .d(input_layer[249]),
      .e(input_layer[381]),
      .f(input_layer[229]),
      .y(Y[1773]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_430 for neuron1774_1
  function_430 neuron1774_1 (
      .a(~input_layer[857]),
      .b(input_layer[306]),
      .c(input_layer[1004]),
      .d(~input_layer[861]),
      .e(input_layer[277]),
      .f(~input_layer[869]),
      .y(Y[1774]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_329 for neuron1775_1
  function_329 neuron1775_1 (
      .a(input_layer[964]),
      .b(~input_layer[452]),
      .c(input_layer[795]),
      .d(~input_layer[382]),
      .e(~input_layer[526]),
      .f(~input_layer[899]),
      .y(Y[1775]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_41 for neuron1776_1
  function_41 neuron1776_1 (
      .a(input_layer[362]),
      .b(input_layer[1279]),
      .c(input_layer[502]),
      .d(~input_layer[659]),
      .e(input_layer[1234]),
      .y(Y[1776]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_363 for neuron1777_1
  function_363 neuron1777_1 (
      .a(~input_layer[1366]),
      .b(~input_layer[648]),
      .c(input_layer[186]),
      .d(~input_layer[1350]),
      .e(input_layer[872]),
      .f(input_layer[742]),
      .y(Y[1777]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1778_1
  function_8 neuron1778_1 (
      .a(input_layer[1493]),
      .b(~input_layer[886]),
      .c(input_layer[732]),
      .d(input_layer[447]),
      .y(Y[1778]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1779_1
  function_299 neuron1779_1 (
      .a(~input_layer[1369]),
      .b(~input_layer[1124]),
      .c(input_layer[201]),
      .d(input_layer[316]),
      .e(~input_layer[370]),
      .y(Y[1779]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron1780_1
  function_75 neuron1780_1 (
      .a(input_layer[514]),
      .b(~input_layer[586]),
      .c(~input_layer[1104]),
      .d(~input_layer[719]),
      .e(input_layer[1496]),
      .y(Y[1780]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_184 for neuron1781_1
  function_184 neuron1781_1 (
      .a(~input_layer[1317]),
      .b(~input_layer[397]),
      .c(input_layer[1325]),
      .d(~input_layer[1017]),
      .e(~input_layer[488]),
      .y(Y[1781]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1782_1
  function_5 neuron1782_1 (
      .a(~input_layer[752]),
      .b(~input_layer[153]),
      .c(~input_layer[613]),
      .d(input_layer[473]),
      .e(~input_layer[1295]),
      .f(input_layer[1407]),
      .y(Y[1782]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1783_1
  function_186 neuron1783_1 (
      .a(~input_layer[496]),
      .b(input_layer[1432]),
      .c(input_layer[1428]),
      .d(~input_layer[594]),
      .y(Y[1783]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1784_1
  function_16 neuron1784_1 (
      .a(~input_layer[580]),
      .b(input_layer[734]),
      .y(Y[1784]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1785_1
  function_67 neuron1785_1 (
      .a(~input_layer[209]),
      .b(~input_layer[182]),
      .c(input_layer[1446]),
      .d(~input_layer[80]),
      .e(~input_layer[374]),
      .y(Y[1785]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron1786_1
  function_290 neuron1786_1 (
      .a(~input_layer[499]),
      .b(~input_layer[1316]),
      .c(~input_layer[1130]),
      .d(input_layer[566]),
      .e(input_layer[1413]),
      .f(input_layer[1233]),
      .y(Y[1786]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron1787_1
  function_175 neuron1787_1 (
      .a(input_layer[318]),
      .b(input_layer[387]),
      .c(input_layer[186]),
      .d(input_layer[748]),
      .e(~input_layer[935]),
      .f(~input_layer[394]),
      .y(Y[1787]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_431 for neuron1788_1
  function_431 neuron1788_1 (
      .a(input_layer[441]),
      .b(~input_layer[190]),
      .c(input_layer[493]),
      .d(input_layer[328]),
      .e(input_layer[743]),
      .f(input_layer[1310]),
      .y(Y[1788]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_346 for neuron1789_1
  function_346 neuron1789_1 (
      .a(~input_layer[1077]),
      .b(input_layer[679]),
      .c(input_layer[717]),
      .d(~input_layer[1292]),
      .e(input_layer[567]),
      .f(input_layer[280]),
      .y(Y[1789]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1790_1
  function_31 neuron1790_1 (
      .a(~input_layer[758]),
      .b(input_layer[774]),
      .c(input_layer[1141]),
      .d(input_layer[527]),
      .y(Y[1790]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron1791_1
  function_84 neuron1791_1 (
      .a(~input_layer[942]),
      .b(input_layer[364]),
      .c(~input_layer[987]),
      .d(~input_layer[98]),
      .e(input_layer[1472]),
      .y(Y[1791]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1792_1
  function_35 neuron1792_1 (
      .a(~input_layer[553]),
      .b(~input_layer[1077]),
      .c(input_layer[708]),
      .d(~input_layer[956]),
      .e(~input_layer[1551]),
      .y(Y[1792]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_432 for neuron1793_1
  function_432 neuron1793_1 (
      .a(~input_layer[798]),
      .b(input_layer[991]),
      .c(~input_layer[1388]),
      .d(input_layer[1303]),
      .e(~input_layer[531]),
      .f(input_layer[96]),
      .y(Y[1793]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1794_1
  function_19 neuron1794_1 (
      .a(~input_layer[1314]),
      .b(~input_layer[613]),
      .c(~input_layer[1252]),
      .d(~input_layer[642]),
      .y(Y[1794]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1795_1
  function_30 neuron1795_1 (
      .a(~input_layer[889]),
      .b(input_layer[235]),
      .c(input_layer[317]),
      .d(~input_layer[1047]),
      .y(Y[1795]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_378 for neuron1796_1
  function_378 neuron1796_1 (
      .a(input_layer[535]),
      .b(~input_layer[1249]),
      .c(input_layer[459]),
      .d(input_layer[471]),
      .e(~input_layer[1284]),
      .f(~input_layer[27]),
      .y(Y[1796]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_314 for neuron1797_1
  function_314 neuron1797_1 (
      .a(input_layer[307]),
      .b(~input_layer[415]),
      .c(~input_layer[576]),
      .d(input_layer[269]),
      .e(~input_layer[578]),
      .y(Y[1797]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_433 for neuron1798_1
  function_433 neuron1798_1 (
      .a(~input_layer[1374]),
      .b(input_layer[146]),
      .c(~input_layer[903]),
      .d(~input_layer[1494]),
      .e(~input_layer[1523]),
      .y(Y[1798]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_434 for neuron1799_1
  function_434 neuron1799_1 (
      .a(input_layer[590]),
      .b(input_layer[517]),
      .c(~input_layer[93]),
      .d(~input_layer[435]),
      .e(input_layer[984]),
      .f(~input_layer[1452]),
      .y(Y[1799]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron1800_1
  function_57 neuron1800_1 (
      .a(input_layer[358]),
      .b(input_layer[989]),
      .c(~input_layer[829]),
      .d(~input_layer[179]),
      .e(input_layer[362]),
      .f(~input_layer[126]),
      .y(Y[1800]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_435 for neuron1801_1
  function_435 neuron1801_1 (
      .a(~input_layer[1416]),
      .b(~input_layer[695]),
      .c(~input_layer[148]),
      .d(input_layer[890]),
      .e(~input_layer[1408]),
      .f(~input_layer[1258]),
      .y(Y[1801]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron1802_1
  function_175 neuron1802_1 (
      .a(input_layer[291]),
      .b(input_layer[933]),
      .c(~input_layer[546]),
      .d(input_layer[444]),
      .e(~input_layer[587]),
      .f(input_layer[955]),
      .y(Y[1802]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_436 for neuron1803_1
  function_436 neuron1803_1 (
      .a(~input_layer[885]),
      .b(~input_layer[1032]),
      .c(~input_layer[1096]),
      .d(input_layer[599]),
      .e(input_layer[600]),
      .f(input_layer[575]),
      .y(Y[1803]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_437 for neuron1804_1
  function_437 neuron1804_1 (
      .a(input_layer[610]),
      .b(~input_layer[586]),
      .c(input_layer[797]),
      .d(~input_layer[884]),
      .e(input_layer[1041]),
      .f(~input_layer[727]),
      .y(Y[1804]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1805_1
  function_27 neuron1805_1 (
      .a(~input_layer[965]),
      .b(input_layer[1359]),
      .c(~input_layer[554]),
      .y(Y[1805]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1806_1
  function_48 neuron1806_1 (
      .a(input_layer[1483]),
      .b(input_layer[702]),
      .c(input_layer[142]),
      .d(~input_layer[598]),
      .e(input_layer[1086]),
      .y(Y[1806]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_438 for neuron1807_1
  function_438 neuron1807_1 (
      .a(~input_layer[694]),
      .b(input_layer[306]),
      .c(input_layer[1552]),
      .d(~input_layer[1271]),
      .e(input_layer[1465]),
      .f(~input_layer[1193]),
      .y(Y[1807]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_129 for neuron1808_1
  function_129 neuron1808_1 (
      .a(~input_layer[699]),
      .b(input_layer[958]),
      .c(input_layer[1467]),
      .d(input_layer[1202]),
      .e(~input_layer[435]),
      .f(~input_layer[1386]),
      .y(Y[1808]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1809_1
  function_12 neuron1809_1 (
      .a(~input_layer[1423]),
      .b(input_layer[1053]),
      .c(input_layer[332]),
      .y(Y[1809]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron1810_1
  function_74 neuron1810_1 (
      .a(~input_layer[831]),
      .b(~input_layer[210]),
      .c(input_layer[708]),
      .d(~input_layer[890]),
      .e(input_layer[354]),
      .f(input_layer[724]),
      .y(Y[1810]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron1811_1
  function_74 neuron1811_1 (
      .a(~input_layer[1473]),
      .b(input_layer[1028]),
      .c(~input_layer[262]),
      .d(input_layer[307]),
      .e(input_layer[1270]),
      .f(~input_layer[1121]),
      .y(Y[1811]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1812] = 1'b1;

  // instantiate function_39 for neuron1813_1
  function_39 neuron1813_1 (
      .a(~input_layer[313]),
      .b(input_layer[1430]),
      .c(~input_layer[800]),
      .y(Y[1813]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_349 for neuron1814_1
  function_349 neuron1814_1 (
      .a(input_layer[566]),
      .b(~input_layer[968]),
      .c(~input_layer[863]),
      .d(input_layer[831]),
      .e(~input_layer[708]),
      .y(Y[1814]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1815_1
  function_3 neuron1815_1 (
      .a(~input_layer[606]),
      .b(~input_layer[830]),
      .c(~input_layer[493]),
      .d(input_layer[652]),
      .y(Y[1815]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1816_1
  function_95 neuron1816_1 (
      .a(input_layer[328]),
      .b(input_layer[1391]),
      .c(~input_layer[1470]),
      .d(~input_layer[737]),
      .y(Y[1816]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron1817_1
  function_61 neuron1817_1 (
      .a(~input_layer[501]),
      .b(input_layer[1107]),
      .c(~input_layer[140]),
      .d(input_layer[778]),
      .e(input_layer[1127]),
      .f(input_layer[1346]),
      .y(Y[1817]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_41 for neuron1818_1
  function_41 neuron1818_1 (
      .a(input_layer[739]),
      .b(input_layer[1364]),
      .c(input_layer[127]),
      .d(input_layer[1556]),
      .e(~input_layer[165]),
      .y(Y[1818]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1819_1
  function_8 neuron1819_1 (
      .a(input_layer[1496]),
      .b(~input_layer[690]),
      .c(input_layer[956]),
      .d(input_layer[1150]),
      .y(Y[1819]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_102 for neuron1820_1
  function_102 neuron1820_1 (
      .a(~input_layer[862]),
      .b(~input_layer[806]),
      .c(~input_layer[363]),
      .d(~input_layer[159]),
      .e(input_layer[602]),
      .f(~input_layer[740]),
      .y(Y[1820]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1821_1
  function_29 neuron1821_1 (
      .a(~input_layer[1084]),
      .b(~input_layer[1085]),
      .y(Y[1821]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1822_1
  function_12 neuron1822_1 (
      .a(~input_layer[437]),
      .b(input_layer[71]),
      .c(input_layer[1339]),
      .y(Y[1822]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1823_1
  function_48 neuron1823_1 (
      .a(input_layer[187]),
      .b(input_layer[134]),
      .c(~input_layer[797]),
      .d(input_layer[97]),
      .e(input_layer[121]),
      .y(Y[1823]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1824_1
  function_26 neuron1824_1 (
      .a(~input_layer[930]),
      .y(Y[1824]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1825_1
  function_106 neuron1825_1 (
      .a(~input_layer[612]),
      .b(input_layer[1103]),
      .c(input_layer[257]),
      .d(input_layer[461]),
      .y(Y[1825]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1826_1
  function_29 neuron1826_1 (
      .a(~input_layer[497]),
      .b(~input_layer[1366]),
      .y(Y[1826]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1827_1
  function_29 neuron1827_1 (
      .a(input_layer[1488]),
      .b(~input_layer[1183]),
      .y(Y[1827]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron1828_1
  function_13 neuron1828_1 (
      .a(input_layer[1216]),
      .b(~input_layer[151]),
      .c(~input_layer[473]),
      .d(~input_layer[1256]),
      .y(Y[1828]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1829_1
  function_16 neuron1829_1 (
      .a(input_layer[926]),
      .b(input_layer[1540]),
      .y(Y[1829]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1830_1
  function_44 neuron1830_1 (
      .a(~input_layer[439]),
      .b(input_layer[598]),
      .c(input_layer[232]),
      .d(~input_layer[1314]),
      .e(~input_layer[305]),
      .y(Y[1830]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_163 for neuron1831_1
  function_163 neuron1831_1 (
      .a(input_layer[648]),
      .b(input_layer[1013]),
      .c(input_layer[412]),
      .d(~input_layer[219]),
      .e(input_layer[276]),
      .y(Y[1831]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1832_1
  function_148 neuron1832_1 (
      .a(input_layer[1472]),
      .b(input_layer[1128]),
      .c(~input_layer[361]),
      .d(~input_layer[1252]),
      .e(input_layer[324]),
      .f(~input_layer[1250]),
      .y(Y[1832]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1833_1
  function_67 neuron1833_1 (
      .a(~input_layer[1147]),
      .b(~input_layer[1061]),
      .c(~input_layer[1501]),
      .d(input_layer[543]),
      .e(~input_layer[619]),
      .y(Y[1833]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1834_1
  function_299 neuron1834_1 (
      .a(input_layer[918]),
      .b(~input_layer[949]),
      .c(~input_layer[78]),
      .d(~input_layer[580]),
      .e(input_layer[1313]),
      .y(Y[1834]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron1835_1
  function_195 neuron1835_1 (
      .a(input_layer[489]),
      .b(input_layer[848]),
      .c(~input_layer[861]),
      .d(input_layer[1251]),
      .e(~input_layer[243]),
      .y(Y[1835]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1836_1
  function_8 neuron1836_1 (
      .a(input_layer[1132]),
      .b(~input_layer[800]),
      .c(input_layer[835]),
      .d(input_layer[234]),
      .y(Y[1836]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_304 for neuron1837_1
  function_304 neuron1837_1 (
      .a(~input_layer[921]),
      .b(~input_layer[1379]),
      .c(input_layer[507]),
      .d(~input_layer[815]),
      .e(~input_layer[367]),
      .f(input_layer[617]),
      .y(Y[1837]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1838_1
  function_47 neuron1838_1 (
      .a(input_layer[1490]),
      .b(input_layer[514]),
      .c(input_layer[316]),
      .d(~input_layer[492]),
      .e(~input_layer[551]),
      .y(Y[1838]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1839_1
  function_26 neuron1839_1 (
      .a(input_layer[491]),
      .y(Y[1839]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1840_1
  function_128 neuron1840_1 (
      .a(~input_layer[974]),
      .b(~input_layer[924]),
      .c(~input_layer[981]),
      .d(input_layer[777]),
      .y(Y[1840]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1841_1
  function_35 neuron1841_1 (
      .a(~input_layer[681]),
      .b(~input_layer[1495]),
      .c(input_layer[253]),
      .d(~input_layer[270]),
      .e(input_layer[347]),
      .y(Y[1841]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_142 for neuron1842_1
  function_142 neuron1842_1 (
      .a(~input_layer[1263]),
      .b(~input_layer[1435]),
      .c(~input_layer[1165]),
      .d(input_layer[232]),
      .e(input_layer[1332]),
      .f(input_layer[1216]),
      .y(Y[1842]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_439 for neuron1843_1
  function_439 neuron1843_1 (
      .a(input_layer[1493]),
      .b(~input_layer[359]),
      .c(input_layer[271]),
      .d(~input_layer[1184]),
      .e(input_layer[530]),
      .f(input_layer[266]),
      .y(Y[1843]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1844_1
  function_8 neuron1844_1 (
      .a(input_layer[586]),
      .b(input_layer[718]),
      .c(~input_layer[1077]),
      .d(~input_layer[186]),
      .y(Y[1844]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1845_1
  function_298 neuron1845_1 (
      .a(~input_layer[145]),
      .b(~input_layer[1199]),
      .c(~input_layer[1010]),
      .d(~input_layer[1397]),
      .e(~input_layer[1394]),
      .f(~input_layer[1565]),
      .y(Y[1845]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron1846_1
  function_241 neuron1846_1 (
      .a(input_layer[852]),
      .b(input_layer[1225]),
      .c(input_layer[1443]),
      .d(input_layer[902]),
      .e(input_layer[473]),
      .f(input_layer[287]),
      .y(Y[1846]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron1847_1
  function_303 neuron1847_1 (
      .a(input_layer[552]),
      .b(input_layer[136]),
      .c(~input_layer[1491]),
      .d(input_layer[1149]),
      .e(input_layer[1267]),
      .f(input_layer[1457]),
      .y(Y[1847]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_417 for neuron1848_1
  function_417 neuron1848_1 (
      .a(~input_layer[432]),
      .b(~input_layer[1433]),
      .c(input_layer[248]),
      .d(~input_layer[633]),
      .e(input_layer[1540]),
      .f(~input_layer[1448]),
      .y(Y[1848]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_222 for neuron1849_1
  function_222 neuron1849_1 (
      .a(input_layer[569]),
      .b(~input_layer[828]),
      .c(input_layer[1276]),
      .d(~input_layer[72]),
      .e(input_layer[19]),
      .f(input_layer[1346]),
      .y(Y[1849]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron1850_1
  function_242 neuron1850_1 (
      .a(input_layer[705]),
      .b(input_layer[1383]),
      .c(input_layer[1327]),
      .d(~input_layer[1103]),
      .e(input_layer[1359]),
      .f(input_layer[730]),
      .y(Y[1850]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1851_1
  function_47 neuron1851_1 (
      .a(input_layer[821]),
      .b(input_layer[139]),
      .c(input_layer[892]),
      .d(input_layer[975]),
      .e(input_layer[276]),
      .y(Y[1851]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron1852_1
  function_6 neuron1852_1 (
      .a(input_layer[368]),
      .b(~input_layer[1449]),
      .c(~input_layer[967]),
      .d(~input_layer[1340]),
      .e(~input_layer[585]),
      .f(input_layer[328]),
      .y(Y[1852]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_440 for neuron1853_1
  function_440 neuron1853_1 (
      .a(~input_layer[246]),
      .b(input_layer[1000]),
      .c(~input_layer[515]),
      .d(~input_layer[123]),
      .e(~input_layer[33]),
      .f(~input_layer[337]),
      .y(Y[1853]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1854_1
  function_16 neuron1854_1 (
      .a(input_layer[579]),
      .b(input_layer[830]),
      .y(Y[1854]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_441 for neuron1855_1
  function_441 neuron1855_1 (
      .a(~input_layer[314]),
      .b(input_layer[1384]),
      .c(~input_layer[461]),
      .d(~input_layer[129]),
      .e(input_layer[707]),
      .f(input_layer[1497]),
      .y(Y[1855]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1856_1
  function_120 neuron1856_1 (
      .a(~input_layer[868]),
      .b(input_layer[87]),
      .c(input_layer[791]),
      .d(input_layer[773]),
      .e(~input_layer[1078]),
      .y(Y[1856]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1857_1
  function_89 neuron1857_1 (
      .a(input_layer[536]),
      .b(~input_layer[885]),
      .c(input_layer[1077]),
      .d(~input_layer[87]),
      .e(input_layer[1349]),
      .y(Y[1857]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_151 for neuron1858_1
  function_151 neuron1858_1 (
      .a(~input_layer[914]),
      .b(input_layer[1350]),
      .c(~input_layer[83]),
      .d(input_layer[1194]),
      .e(~input_layer[1395]),
      .f(~input_layer[1271]),
      .y(Y[1858]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1859_1
  function_42 neuron1859_1 (
      .a(input_layer[877]),
      .b(input_layer[521]),
      .c(input_layer[611]),
      .d(input_layer[891]),
      .y(Y[1859]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1860_1
  function_3 neuron1860_1 (
      .a(~input_layer[1184]),
      .b(~input_layer[356]),
      .c(~input_layer[779]),
      .d(input_layer[814]),
      .y(Y[1860]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1861_1
  function_72 neuron1861_1 (
      .a(input_layer[564]),
      .b(~input_layer[419]),
      .c(~input_layer[365]),
      .d(~input_layer[1488]),
      .e(input_layer[955]),
      .y(Y[1861]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1862_1
  function_17 neuron1862_1 (
      .a(input_layer[1131]),
      .b(input_layer[537]),
      .c(input_layer[1257]),
      .y(Y[1862]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron1863_1
  function_155 neuron1863_1 (
      .a(~input_layer[830]),
      .b(~input_layer[1016]),
      .c(~input_layer[533]),
      .d(~input_layer[721]),
      .e(input_layer[743]),
      .f(~input_layer[75]),
      .y(Y[1863]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1864_1
  function_48 neuron1864_1 (
      .a(input_layer[352]),
      .b(input_layer[602]),
      .c(~input_layer[702]),
      .d(input_layer[545]),
      .e(input_layer[809]),
      .y(Y[1864]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_279 for neuron1865_1
  function_279 neuron1865_1 (
      .a(input_layer[1419]),
      .b(~input_layer[914]),
      .c(~input_layer[943]),
      .d(input_layer[1447]),
      .e(~input_layer[79]),
      .y(Y[1865]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1866] = 1'b0;

  // instantiate function_67 for neuron1867_1
  function_67 neuron1867_1 (
      .a(~input_layer[771]),
      .b(input_layer[408]),
      .c(~input_layer[556]),
      .d(~input_layer[681]),
      .e(~input_layer[886]),
      .y(Y[1867]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1868_1
  function_169 neuron1868_1 (
      .a(~input_layer[365]),
      .b(~input_layer[1276]),
      .c(input_layer[1113]),
      .d(input_layer[64]),
      .e(~input_layer[7]),
      .f(input_layer[3]),
      .y(Y[1868]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1869_1
  function_42 neuron1869_1 (
      .a(input_layer[190]),
      .b(~input_layer[921]),
      .c(input_layer[1468]),
      .d(input_layer[401]),
      .y(Y[1869]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_51 for neuron1870_1
  function_51 neuron1870_1 (
      .a(input_layer[752]),
      .b(~input_layer[1034]),
      .c(~input_layer[524]),
      .d(input_layer[489]),
      .e(~input_layer[832]),
      .f(~input_layer[1289]),
      .y(Y[1870]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_442 for neuron1871_1
  function_442 neuron1871_1 (
      .a(input_layer[188]),
      .b(~input_layer[852]),
      .c(~input_layer[707]),
      .d(~input_layer[793]),
      .e(input_layer[734]),
      .f(~input_layer[162]),
      .y(Y[1871]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1872_1
  function_0 neuron1872_1 (
      .a(~input_layer[998]),
      .b(~input_layer[1117]),
      .c(~input_layer[1229]),
      .d(~input_layer[1008]),
      .e(input_layer[1346]),
      .y(Y[1872]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1873_1
  function_17 neuron1873_1 (
      .a(input_layer[753]),
      .b(input_layer[1182]),
      .c(input_layer[332]),
      .y(Y[1873]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_58 for neuron1874_1
  function_58 neuron1874_1 (
      .a(input_layer[719]),
      .b(~input_layer[634]),
      .c(input_layer[1300]),
      .d(input_layer[1205]),
      .e(input_layer[1073]),
      .f(~input_layer[684]),
      .y(Y[1874]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1875_1
  function_27 neuron1875_1 (
      .a(~input_layer[1167]),
      .b(~input_layer[252]),
      .c(~input_layer[991]),
      .y(Y[1875]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1876_1
  function_167 neuron1876_1 (
      .a(input_layer[827]),
      .b(input_layer[879]),
      .c(input_layer[697]),
      .d(~input_layer[867]),
      .e(input_layer[90]),
      .y(Y[1876]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_443 for neuron1877_1
  function_443 neuron1877_1 (
      .a(input_layer[808]),
      .b(~input_layer[775]),
      .c(input_layer[88]),
      .d(input_layer[1357]),
      .e(input_layer[1292]),
      .f(input_layer[620]),
      .y(Y[1877]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_238 for neuron1878_1
  function_238 neuron1878_1 (
      .a(input_layer[1073]),
      .b(~input_layer[197]),
      .c(~input_layer[92]),
      .d(input_layer[353]),
      .e(~input_layer[177]),
      .y(Y[1878]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_444 for neuron1879_1
  function_444 neuron1879_1 (
      .a(input_layer[579]),
      .b(~input_layer[1113]),
      .c(input_layer[1443]),
      .d(input_layer[437]),
      .e(~input_layer[1116]),
      .f(~input_layer[1422]),
      .y(Y[1879]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_445 for neuron1880_1
  function_445 neuron1880_1 (
      .a(input_layer[1274]),
      .b(~input_layer[768]),
      .c(~input_layer[212]),
      .d(input_layer[707]),
      .e(input_layer[1173]),
      .f(~input_layer[1211]),
      .y(Y[1880]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1881_1
  function_135 neuron1881_1 (
      .a(input_layer[1215]),
      .b(~input_layer[1543]),
      .c(~input_layer[531]),
      .d(input_layer[355]),
      .e(input_layer[831]),
      .y(Y[1881]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1882_1
  function_47 neuron1882_1 (
      .a(input_layer[425]),
      .b(input_layer[374]),
      .c(input_layer[1280]),
      .d(~input_layer[1151]),
      .e(input_layer[1263]),
      .y(Y[1882]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1883_1
  function_27 neuron1883_1 (
      .a(~input_layer[767]),
      .b(~input_layer[150]),
      .c(input_layer[491]),
      .y(Y[1883]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1884_1
  function_35 neuron1884_1 (
      .a(~input_layer[185]),
      .b(input_layer[917]),
      .c(~input_layer[1217]),
      .d(input_layer[969]),
      .e(~input_layer[640]),
      .y(Y[1884]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1885_1
  function_92 neuron1885_1 (
      .a(input_layer[858]),
      .b(input_layer[1124]),
      .c(input_layer[938]),
      .d(input_layer[820]),
      .e(input_layer[741]),
      .f(input_layer[1195]),
      .y(Y[1885]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1886_1
  function_100 neuron1886_1 (
      .a(~input_layer[477]),
      .b(~input_layer[1237]),
      .c(~input_layer[781]),
      .d(~input_layer[1011]),
      .e(input_layer[295]),
      .f(~input_layer[569]),
      .y(Y[1886]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1887_1
  function_0 neuron1887_1 (
      .a(~input_layer[1418]),
      .b(~input_layer[474]),
      .c(~input_layer[933]),
      .d(~input_layer[1326]),
      .e(~input_layer[488]),
      .y(Y[1887]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1888_1
  function_42 neuron1888_1 (
      .a(input_layer[213]),
      .b(input_layer[184]),
      .c(input_layer[1203]),
      .d(input_layer[80]),
      .y(Y[1888]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1889_1
  function_39 neuron1889_1 (
      .a(~input_layer[209]),
      .b(input_layer[1423]),
      .c(input_layer[482]),
      .y(Y[1889]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1890_1
  function_24 neuron1890_1 (
      .a(~input_layer[1034]),
      .b(input_layer[1262]),
      .c(~input_layer[606]),
      .y(Y[1890]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_446 for neuron1891_1
  function_446 neuron1891_1 (
      .a(input_layer[1107]),
      .b(~input_layer[792]),
      .c(~input_layer[29]),
      .d(~input_layer[17]),
      .e(input_layer[617]),
      .f(~input_layer[1015]),
      .y(Y[1891]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_447 for neuron1892_1
  function_447 neuron1892_1 (
      .a(~input_layer[1473]),
      .b(input_layer[183]),
      .c(input_layer[1192]),
      .d(~input_layer[1489]),
      .e(input_layer[426]),
      .f(~input_layer[572]),
      .y(Y[1892]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1893_1
  function_8 neuron1893_1 (
      .a(input_layer[1226]),
      .b(input_layer[987]),
      .c(~input_layer[850]),
      .d(input_layer[1095]),
      .y(Y[1893]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1894_1
  function_0 neuron1894_1 (
      .a(~input_layer[1050]),
      .b(input_layer[1495]),
      .c(~input_layer[89]),
      .d(~input_layer[901]),
      .e(~input_layer[413]),
      .y(Y[1894]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1895_1
  function_17 neuron1895_1 (
      .a(input_layer[656]),
      .b(input_layer[309]),
      .c(input_layer[471]),
      .y(Y[1895]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1896_1
  function_89 neuron1896_1 (
      .a(input_layer[354]),
      .b(~input_layer[876]),
      .c(~input_layer[1432]),
      .d(input_layer[1525]),
      .e(input_layer[161]),
      .y(Y[1896]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1897_1
  function_27 neuron1897_1 (
      .a(~input_layer[829]),
      .b(~input_layer[777]),
      .c(~input_layer[750]),
      .y(Y[1897]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1898_1
  function_154 neuron1898_1 (
      .a(~input_layer[640]),
      .b(~input_layer[499]),
      .c(input_layer[910]),
      .d(~input_layer[1549]),
      .e(input_layer[1234]),
      .f(input_layer[834]),
      .y(Y[1898]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_108 for neuron1899_1
  function_108 neuron1899_1 (
      .a(input_layer[1299]),
      .b(input_layer[1250]),
      .c(input_layer[1315]),
      .d(input_layer[1265]),
      .e(~input_layer[807]),
      .f(input_layer[1217]),
      .y(Y[1899]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1900_1
  function_90 neuron1900_1 (
      .a(~input_layer[918]),
      .b(~input_layer[861]),
      .c(~input_layer[1332]),
      .d(input_layer[1039]),
      .e(~input_layer[608]),
      .y(Y[1900]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1901_1
  function_27 neuron1901_1 (
      .a(input_layer[1032]),
      .b(~input_layer[1484]),
      .c(~input_layer[627]),
      .y(Y[1901]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron1902_1
  function_286 neuron1902_1 (
      .a(input_layer[761]),
      .b(~input_layer[372]),
      .c(~input_layer[360]),
      .d(~input_layer[94]),
      .e(~input_layer[229]),
      .y(Y[1902]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1903_1
  function_271 neuron1903_1 (
      .a(input_layer[1188]),
      .b(input_layer[1185]),
      .c(input_layer[241]),
      .d(~input_layer[1323]),
      .e(~input_layer[697]),
      .y(Y[1903]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_448 for neuron1904_1
  function_448 neuron1904_1 (
      .a(~input_layer[304]),
      .b(input_layer[1496]),
      .c(~input_layer[394]),
      .d(input_layer[160]),
      .e(~input_layer[785]),
      .y(Y[1904]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1905_1
  function_1 neuron1905_1 (
      .a(input_layer[138]),
      .b(~input_layer[1272]),
      .c(~input_layer[318]),
      .d(~input_layer[432]),
      .y(Y[1905]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron1906_1
  function_192 neuron1906_1 (
      .a(~input_layer[981]),
      .b(input_layer[717]),
      .c(input_layer[75]),
      .d(~input_layer[737]),
      .e(input_layer[428]),
      .f(input_layer[1349]),
      .y(Y[1906]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1907_1
  function_55 neuron1907_1 (
      .a(~input_layer[938]),
      .b(input_layer[651]),
      .c(~input_layer[1133]),
      .d(~input_layer[679]),
      .e(~input_layer[779]),
      .y(Y[1907]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1908_1
  function_3 neuron1908_1 (
      .a(~input_layer[407]),
      .b(~input_layer[875]),
      .c(~input_layer[941]),
      .d(~input_layer[724]),
      .y(Y[1908]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_449 for neuron1909_1
  function_449 neuron1909_1 (
      .a(input_layer[1439]),
      .b(input_layer[1489]),
      .c(input_layer[764]),
      .d(~input_layer[344]),
      .e(~input_layer[677]),
      .y(Y[1909]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_354 for neuron1910_1
  function_354 neuron1910_1 (
      .a(input_layer[964]),
      .b(~input_layer[76]),
      .c(~input_layer[308]),
      .d(~input_layer[24]),
      .e(input_layer[1455]),
      .f(~input_layer[50]),
      .y(Y[1910]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_363 for neuron1911_1
  function_363 neuron1911_1 (
      .a(~input_layer[609]),
      .b(input_layer[1236]),
      .c(input_layer[126]),
      .d(~input_layer[1410]),
      .e(input_layer[1404]),
      .f(~input_layer[334]),
      .y(Y[1911]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1912_1
  function_7 neuron1912_1 (
      .a(~input_layer[534]),
      .b(input_layer[804]),
      .c(~input_layer[1208]),
      .d(input_layer[1063]),
      .y(Y[1912]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_450 for neuron1913_1
  function_450 neuron1913_1 (
      .a(~input_layer[833]),
      .b(input_layer[445]),
      .c(input_layer[1252]),
      .d(input_layer[1115]),
      .e(input_layer[1137]),
      .f(~input_layer[1211]),
      .y(Y[1913]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1914_1
  function_19 neuron1914_1 (
      .a(~input_layer[607]),
      .b(input_layer[1039]),
      .c(~input_layer[489]),
      .d(~input_layer[99]),
      .y(Y[1914]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron1915_1
  function_78 neuron1915_1 (
      .a(~input_layer[479]),
      .b(~input_layer[1296]),
      .c(~input_layer[1533]),
      .d(input_layer[929]),
      .e(~input_layer[548]),
      .f(input_layer[920]),
      .y(Y[1915]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron1916_1
  function_59 neuron1916_1 (
      .a(~input_layer[757]),
      .b(input_layer[405]),
      .c(input_layer[1223]),
      .d(input_layer[275]),
      .e(input_layer[742]),
      .f(~input_layer[75]),
      .y(Y[1916]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron1917_1
  function_221 neuron1917_1 (
      .a(input_layer[415]),
      .b(~input_layer[871]),
      .c(input_layer[714]),
      .d(input_layer[1431]),
      .e(~input_layer[459]),
      .f(input_layer[1554]),
      .y(Y[1917]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1918_1
  function_181 neuron1918_1 (
      .a(input_layer[1375]),
      .b(~input_layer[1087]),
      .c(~input_layer[1488]),
      .d(~input_layer[1553]),
      .e(input_layer[954]),
      .y(Y[1918]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1919_1
  function_24 neuron1919_1 (
      .a(~input_layer[1252]),
      .b(input_layer[264]),
      .c(~input_layer[1218]),
      .y(Y[1919]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_451 for neuron1920_1
  function_451 neuron1920_1 (
      .a(~input_layer[705]),
      .b(~input_layer[572]),
      .c(input_layer[381]),
      .d(input_layer[531]),
      .e(~input_layer[836]),
      .f(~input_layer[606]),
      .y(Y[1920]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1921_1
  function_24 neuron1921_1 (
      .a(~input_layer[581]),
      .b(input_layer[596]),
      .c(input_layer[1322]),
      .y(Y[1921]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1922] = 1'b1;

  // instantiate function_291 for neuron1923_1
  function_291 neuron1923_1 (
      .a(input_layer[972]),
      .b(input_layer[968]),
      .c(~input_layer[623]),
      .d(input_layer[865]),
      .e(input_layer[160]),
      .y(Y[1923]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1924_1
  function_3 neuron1924_1 (
      .a(~input_layer[884]),
      .b(~input_layer[1182]),
      .c(~input_layer[704]),
      .d(~input_layer[835]),
      .y(Y[1924]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1925_1
  function_27 neuron1925_1 (
      .a(~input_layer[1424]),
      .b(~input_layer[1283]),
      .c(input_layer[864]),
      .y(Y[1925]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1926_1
  function_17 neuron1926_1 (
      .a(input_layer[871]),
      .b(input_layer[202]),
      .c(input_layer[327]),
      .y(Y[1926]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1927_1
  function_7 neuron1927_1 (
      .a(input_layer[1475]),
      .b(~input_layer[238]),
      .c(input_layer[707]),
      .d(input_layer[26]),
      .y(Y[1927]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_205 for neuron1928_1
  function_205 neuron1928_1 (
      .a(input_layer[918]),
      .b(~input_layer[1334]),
      .c(input_layer[200]),
      .d(~input_layer[1444]),
      .e(~input_layer[1534]),
      .f(input_layer[27]),
      .y(Y[1928]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1929_1
  function_47 neuron1929_1 (
      .a(input_layer[182]),
      .b(input_layer[81]),
      .c(~input_layer[1084]),
      .d(~input_layer[1260]),
      .e(input_layer[125]),
      .y(Y[1929]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1930_1
  function_87 neuron1930_1 (
      .a(input_layer[1376]),
      .b(~input_layer[993]),
      .c(~input_layer[825]),
      .d(input_layer[452]),
      .e(input_layer[1503]),
      .y(Y[1930]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1931_1
  function_30 neuron1931_1 (
      .a(input_layer[1136]),
      .b(~input_layer[814]),
      .c(~input_layer[1335]),
      .d(input_layer[573]),
      .y(Y[1931]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1932_1
  function_48 neuron1932_1 (
      .a(input_layer[1493]),
      .b(input_layer[1171]),
      .c(input_layer[1217]),
      .d(input_layer[1283]),
      .e(~input_layer[265]),
      .y(Y[1932]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron1933_1
  function_242 neuron1933_1 (
      .a(input_layer[1475]),
      .b(~input_layer[1079]),
      .c(input_layer[541]),
      .d(input_layer[844]),
      .e(input_layer[1063]),
      .f(input_layer[1066]),
      .y(Y[1933]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_412 for neuron1934_1
  function_412 neuron1934_1 (
      .a(input_layer[857]),
      .b(~input_layer[703]),
      .c(input_layer[626]),
      .d(~input_layer[72]),
      .e(input_layer[430]),
      .y(Y[1934]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron1935_1
  function_241 neuron1935_1 (
      .a(input_layer[508]),
      .b(input_layer[1359]),
      .c(~input_layer[1119]),
      .d(input_layer[177]),
      .e(input_layer[7]),
      .f(input_layer[1120]),
      .y(Y[1935]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_452 for neuron1936_1
  function_452 neuron1936_1 (
      .a(input_layer[703]),
      .b(~input_layer[147]),
      .c(~input_layer[444]),
      .d(input_layer[240]),
      .e(~input_layer[432]),
      .f(~input_layer[486]),
      .y(Y[1936]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron1937_1
  function_186 neuron1937_1 (
      .a(~input_layer[1035]),
      .b(input_layer[721]),
      .c(~input_layer[1277]),
      .d(input_layer[577]),
      .y(Y[1937]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1938_1
  function_17 neuron1938_1 (
      .a(input_layer[904]),
      .b(~input_layer[1322]),
      .c(input_layer[1203]),
      .y(Y[1938]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1939_1
  function_4 neuron1939_1 (
      .a(~input_layer[1126]),
      .b(~input_layer[1534]),
      .c(input_layer[594]),
      .d(~input_layer[662]),
      .e(~input_layer[843]),
      .y(Y[1939]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1940_1
  function_24 neuron1940_1 (
      .a(~input_layer[1206]),
      .b(~input_layer[465]),
      .c(input_layer[944]),
      .y(Y[1940]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1941_1
  function_172 neuron1941_1 (
      .a(~input_layer[202]),
      .b(~input_layer[1159]),
      .c(~input_layer[1001]),
      .d(input_layer[870]),
      .e(input_layer[1446]),
      .f(~input_layer[780]),
      .y(Y[1941]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1942_1
  function_299 neuron1942_1 (
      .a(input_layer[347]),
      .b(~input_layer[1442]),
      .c(~input_layer[1263]),
      .d(~input_layer[127]),
      .e(~input_layer[124]),
      .y(Y[1942]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1943_1
  function_146 neuron1943_1 (
      .a(input_layer[247]),
      .b(input_layer[1367]),
      .c(input_layer[555]),
      .d(~input_layer[691]),
      .e(input_layer[943]),
      .f(input_layer[755]),
      .y(Y[1943]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron1944_1
  function_57 neuron1944_1 (
      .a(~input_layer[591]),
      .b(input_layer[1381]),
      .c(input_layer[100]),
      .d(~input_layer[220]),
      .e(input_layer[1513]),
      .f(input_layer[72]),
      .y(Y[1944]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1945_1
  function_91 neuron1945_1 (
      .a(~input_layer[554]),
      .b(input_layer[138]),
      .c(input_layer[251]),
      .d(input_layer[1048]),
      .e(~input_layer[1357]),
      .y(Y[1945]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1946_1
  function_28 neuron1946_1 (
      .a(~input_layer[459]),
      .b(~input_layer[888]),
      .c(~input_layer[91]),
      .d(~input_layer[90]),
      .e(~input_layer[1426]),
      .f(input_layer[1321]),
      .y(Y[1946]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1947_1
  function_31 neuron1947_1 (
      .a(input_layer[428]),
      .b(~input_layer[182]),
      .c(~input_layer[832]),
      .d(input_layer[629]),
      .y(Y[1947]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_220 for neuron1948_1
  function_220 neuron1948_1 (
      .a(~input_layer[923]),
      .b(input_layer[797]),
      .c(input_layer[769]),
      .d(input_layer[1165]),
      .e(input_layer[322]),
      .f(input_layer[1563]),
      .y(Y[1948]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_453 for neuron1949_1
  function_453 neuron1949_1 (
      .a(input_layer[483]),
      .b(input_layer[959]),
      .c(~input_layer[966]),
      .d(~input_layer[796]),
      .e(~input_layer[179]),
      .f(~input_layer[27]),
      .y(Y[1949]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron1950_1
  function_165 neuron1950_1 (
      .a(input_layer[773]),
      .b(~input_layer[1252]),
      .c(~input_layer[1181]),
      .d(input_layer[663]),
      .e(~input_layer[1558]),
      .y(Y[1950]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_206 for neuron1951_1
  function_206 neuron1951_1 (
      .a(~input_layer[467]),
      .b(~input_layer[488]),
      .c(~input_layer[1182]),
      .d(input_layer[1201]),
      .e(~input_layer[1348]),
      .f(input_layer[1555]),
      .y(Y[1951]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1952_1
  function_48 neuron1952_1 (
      .a(input_layer[1239]),
      .b(input_layer[1472]),
      .c(~input_layer[925]),
      .d(input_layer[1535]),
      .e(~input_layer[386]),
      .y(Y[1952]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_151 for neuron1953_1
  function_151 neuron1953_1 (
      .a(input_layer[1030]),
      .b(~input_layer[409]),
      .c(~input_layer[655]),
      .d(~input_layer[232]),
      .e(input_layer[203]),
      .f(~input_layer[1234]),
      .y(Y[1953]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron1954_1
  function_47 neuron1954_1 (
      .a(input_layer[599]),
      .b(input_layer[716]),
      .c(input_layer[774]),
      .d(input_layer[1027]),
      .e(~input_layer[372]),
      .y(Y[1954]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron1955_1
  function_6 neuron1955_1 (
      .a(~input_layer[654]),
      .b(~input_layer[88]),
      .c(~input_layer[295]),
      .d(input_layer[1236]),
      .e(~input_layer[1535]),
      .f(~input_layer[1550]),
      .y(Y[1955]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1956_1
  function_67 neuron1956_1 (
      .a(input_layer[927]),
      .b(~input_layer[1060]),
      .c(~input_layer[1542]),
      .d(~input_layer[1466]),
      .e(~input_layer[452]),
      .y(Y[1956]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1957_1
  function_26 neuron1957_1 (
      .a(input_layer[761]),
      .y(Y[1957]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1958_1
  function_35 neuron1958_1 (
      .a(~input_layer[991]),
      .b(input_layer[706]),
      .c(~input_layer[891]),
      .d(~input_layer[1023]),
      .e(~input_layer[30]),
      .y(Y[1958]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1959_1
  function_26 neuron1959_1 (
      .a(input_layer[1250]),
      .y(Y[1959]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1960_1
  function_123 neuron1960_1 (
      .a(input_layer[976]),
      .b(input_layer[1226]),
      .c(~input_layer[457]),
      .d(~input_layer[674]),
      .y(Y[1960]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1961_1
  function_17 neuron1961_1 (
      .a(input_layer[1216]),
      .b(input_layer[1494]),
      .c(input_layer[1536]),
      .y(Y[1961]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1962_1
  function_92 neuron1962_1 (
      .a(input_layer[141]),
      .b(input_layer[292]),
      .c(~input_layer[472]),
      .d(input_layer[1002]),
      .e(~input_layer[576]),
      .f(input_layer[786]),
      .y(Y[1962]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron1963_1
  function_55 neuron1963_1 (
      .a(~input_layer[1015]),
      .b(~input_layer[1005]),
      .c(~input_layer[1411]),
      .d(input_layer[1038]),
      .e(input_layer[1331]),
      .y(Y[1963]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1964_1
  function_8 neuron1964_1 (
      .a(input_layer[422]),
      .b(input_layer[1059]),
      .c(input_layer[235]),
      .d(input_layer[122]),
      .y(Y[1964]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_454 for neuron1965_1
  function_454 neuron1965_1 (
      .a(~input_layer[580]),
      .b(input_layer[1171]),
      .c(input_layer[905]),
      .d(input_layer[234]),
      .e(~input_layer[549]),
      .f(~input_layer[1391]),
      .y(Y[1965]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron1966_1
  function_271 neuron1966_1 (
      .a(input_layer[313]),
      .b(~input_layer[464]),
      .c(input_layer[1171]),
      .d(~input_layer[628]),
      .e(input_layer[836]),
      .y(Y[1966]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1967_1
  function_1 neuron1967_1 (
      .a(~input_layer[482]),
      .b(~input_layer[1530]),
      .c(input_layer[710]),
      .d(input_layer[1229]),
      .y(Y[1967]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron1968_1
  function_8 neuron1968_1 (
      .a(input_layer[995]),
      .b(~input_layer[370]),
      .c(input_layer[1393]),
      .d(input_layer[845]),
      .y(Y[1968]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron1969_1
  function_121 neuron1969_1 (
      .a(input_layer[775]),
      .b(input_layer[1440]),
      .c(~input_layer[1245]),
      .d(input_layer[922]),
      .e(input_layer[1084]),
      .y(Y[1969]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1970_1
  function_29 neuron1970_1 (
      .a(~input_layer[936]),
      .b(~input_layer[461]),
      .y(Y[1970]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron1971_1
  function_42 neuron1971_1 (
      .a(input_layer[579]),
      .b(input_layer[1270]),
      .c(input_layer[155]),
      .d(input_layer[1051]),
      .y(Y[1971]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1972_1
  function_11 neuron1972_1 (
      .a(input_layer[355]),
      .b(~input_layer[1275]),
      .c(~input_layer[1148]),
      .d(~input_layer[789]),
      .y(Y[1972]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron1973_1
  function_106 neuron1973_1 (
      .a(input_layer[651]),
      .b(~input_layer[807]),
      .c(~input_layer[804]),
      .d(input_layer[877]),
      .y(Y[1973]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1974_1
  function_330 neuron1974_1 (
      .a(~input_layer[1073]),
      .b(~input_layer[1314]),
      .c(input_layer[626]),
      .d(input_layer[618]),
      .e(input_layer[731]),
      .y(Y[1974]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_446 for neuron1975_1
  function_446 neuron1975_1 (
      .a(input_layer[752]),
      .b(input_layer[254]),
      .c(~input_layer[518]),
      .d(input_layer[1377]),
      .e(input_layer[96]),
      .f(~input_layer[228]),
      .y(Y[1975]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron1976_1
  function_27 neuron1976_1 (
      .a(~input_layer[1352]),
      .b(input_layer[303]),
      .c(~input_layer[69]),
      .y(Y[1976]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron1977_1
  function_29 neuron1977_1 (
      .a(~input_layer[429]),
      .b(~input_layer[475]),
      .y(Y[1977]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_455 for neuron1978_1
  function_455 neuron1978_1 (
      .a(~input_layer[1221]),
      .b(input_layer[868]),
      .c(~input_layer[1027]),
      .d(input_layer[1353]),
      .e(~input_layer[430]),
      .f(~input_layer[1071]),
      .y(Y[1978]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_456 for neuron1979_1
  function_456 neuron1979_1 (
      .a(input_layer[1490]),
      .b(~input_layer[911]),
      .c(input_layer[562]),
      .d(input_layer[451]),
      .e(~input_layer[539]),
      .f(input_layer[1328]),
      .y(Y[1979]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1980_1
  function_17 neuron1980_1 (
      .a(input_layer[604]),
      .b(input_layer[1111]),
      .c(input_layer[216]),
      .y(Y[1980]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron1981_1
  function_7 neuron1981_1 (
      .a(input_layer[1434]),
      .b(~input_layer[596]),
      .c(input_layer[1430]),
      .d(~input_layer[177]),
      .y(Y[1981]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_218 for neuron1982_1
  function_218 neuron1982_1 (
      .a(input_layer[205]),
      .b(input_layer[443]),
      .c(~input_layer[1370]),
      .d(~input_layer[743]),
      .e(input_layer[1090]),
      .y(Y[1982]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_251 for neuron1983_1
  function_251 neuron1983_1 (
      .a(input_layer[908]),
      .b(~input_layer[1111]),
      .c(input_layer[309]),
      .d(~input_layer[1079]),
      .e(input_layer[1525]),
      .f(input_layer[129]),
      .y(Y[1983]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_457 for neuron1984_1
  function_457 neuron1984_1 (
      .a(~input_layer[608]),
      .b(input_layer[657]),
      .c(~input_layer[129]),
      .d(input_layer[1334]),
      .e(input_layer[1497]),
      .f(~input_layer[770]),
      .y(Y[1984]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1985_1
  function_87 neuron1985_1 (
      .a(input_layer[1018]),
      .b(input_layer[1137]),
      .c(input_layer[985]),
      .d(~input_layer[400]),
      .e(~input_layer[933]),
      .y(Y[1985]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1986_1
  function_26 neuron1986_1 (
      .a(~input_layer[1042]),
      .y(Y[1986]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1987_1
  function_3 neuron1987_1 (
      .a(~input_layer[152]),
      .b(~input_layer[1247]),
      .c(~input_layer[154]),
      .d(input_layer[708]),
      .y(Y[1987]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1988_1
  function_104 neuron1988_1 (
      .a(~input_layer[932]),
      .b(input_layer[1436]),
      .c(~input_layer[1106]),
      .d(input_layer[712]),
      .e(input_layer[1558]),
      .f(input_layer[896]),
      .y(Y[1988]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron1989_1
  function_97 neuron1989_1 (
      .a(~input_layer[656]),
      .b(~input_layer[235]),
      .c(~input_layer[927]),
      .d(input_layer[333]),
      .e(~input_layer[1390]),
      .y(Y[1989]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_397 for neuron1990_1
  function_397 neuron1990_1 (
      .a(input_layer[1539]),
      .b(~input_layer[1371]),
      .c(~input_layer[549]),
      .d(input_layer[836]),
      .e(~input_layer[865]),
      .y(Y[1990]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1991_1
  function_113 neuron1991_1 (
      .a(input_layer[973]),
      .b(input_layer[682]),
      .c(~input_layer[189]),
      .d(~input_layer[541]),
      .e(input_layer[324]),
      .y(Y[1991]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1992_1
  function_17 neuron1992_1 (
      .a(input_layer[760]),
      .b(input_layer[1431]),
      .c(input_layer[205]),
      .y(Y[1992]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1993_1
  function_135 neuron1993_1 (
      .a(input_layer[539]),
      .b(~input_layer[831]),
      .c(input_layer[679]),
      .d(input_layer[652]),
      .e(~input_layer[982]),
      .y(Y[1993]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron1994_1
  function_46 neuron1994_1 (
      .a(input_layer[1087]),
      .b(input_layer[1059]),
      .c(input_layer[206]),
      .d(~input_layer[1236]),
      .e(~input_layer[462]),
      .y(Y[1994]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_419 for neuron1995_1
  function_419 neuron1995_1 (
      .a(~input_layer[419]),
      .b(input_layer[585]),
      .c(input_layer[856]),
      .d(input_layer[578]),
      .e(input_layer[747]),
      .f(~input_layer[592]),
      .y(Y[1995]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1996_1
  function_31 neuron1996_1 (
      .a(input_layer[190]),
      .b(~input_layer[1423]),
      .c(~input_layer[654]),
      .d(input_layer[917]),
      .y(Y[1996]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron1997_1
  function_156 neuron1997_1 (
      .a(~input_layer[1151]),
      .b(~input_layer[436]),
      .c(~input_layer[1230]),
      .d(input_layer[785]),
      .e(~input_layer[1563]),
      .f(~input_layer[726]),
      .y(Y[1997]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_23 for neuron1998_1
  function_23 neuron1998_1 (
      .a(~input_layer[437]),
      .b(~input_layer[306]),
      .c(input_layer[572]),
      .d(~input_layer[1254]),
      .e(input_layer[1286]),
      .f(~input_layer[956]),
      .y(Y[1998]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron1999_1
  function_195 neuron1999_1 (
      .a(input_layer[638]),
      .b(~input_layer[978]),
      .c(input_layer[854]),
      .d(~input_layer[999]),
      .e(input_layer[1261]),
      .y(Y[1999]),
      .clk(clk),
      .rst(rst)
  );

// total zero consts: 23
// total one  consts: 13
// total instantiations: 1964

  // Warning: Z[0] not driven (layer 3)
  // Warning: Z[1] not driven (layer 3)
  // Warning: Z[2] not driven (layer 3)
  // Warning: Z[3] not driven (layer 3)
  // Warning: Z[4] not driven (layer 3)
  // Warning: Z[5] not driven (layer 3)
  // Warning: Z[6] not driven (layer 3)
  // Warning: Z[7] not driven (layer 3)
  // Warning: Z[8] not driven (layer 3)
  // Warning: Z[9] not driven (layer 3)
  // Warning: Z[10] not driven (layer 3)
  // Warning: Z[11] not driven (layer 3)
  // Warning: Z[12] not driven (layer 3)
  // Warning: Z[13] not driven (layer 3)
  // Warning: Z[14] not driven (layer 3)
  // Warning: Z[15] not driven (layer 3)
  // Warning: Z[16] not driven (layer 3)
  // Warning: Z[17] not driven (layer 3)
  // Warning: Z[18] not driven (layer 3)
  // Warning: Z[19] not driven (layer 3)
  // Warning: Z[20] not driven (layer 3)
  // Warning: Z[21] not driven (layer 3)
  // Warning: Z[22] not driven (layer 3)
  // Warning: Z[23] not driven (layer 3)
  // Warning: Z[24] not driven (layer 3)
  // Warning: Z[25] not driven (layer 3)
  // Warning: Z[26] not driven (layer 3)
  // Warning: Z[27] not driven (layer 3)
  // Warning: Z[28] not driven (layer 3)
  // Warning: Z[29] not driven (layer 3)
  // Warning: Z[30] not driven (layer 3)
  // Warning: Z[31] not driven (layer 3)
  // Warning: Z[32] not driven (layer 3)
  // Warning: Z[33] not driven (layer 3)
  // Warning: Z[34] not driven (layer 3)
  // Warning: Z[35] not driven (layer 3)
  // Warning: Z[36] not driven (layer 3)
  // Warning: Z[37] not driven (layer 3)
  // Warning: Z[38] not driven (layer 3)
  // Warning: Z[39] not driven (layer 3)
  // Warning: Z[40] not driven (layer 3)
  // Warning: Z[41] not driven (layer 3)
  // Warning: Z[42] not driven (layer 3)
  // Warning: Z[43] not driven (layer 3)
  // Warning: Z[44] not driven (layer 3)
  // Warning: Z[45] not driven (layer 3)
  // Warning: Z[46] not driven (layer 3)
  // Warning: Z[47] not driven (layer 3)
  // Warning: Z[48] not driven (layer 3)
  // Warning: Z[49] not driven (layer 3)
  // Warning: Z[50] not driven (layer 3)
  // Warning: Z[51] not driven (layer 3)
  // Warning: Z[52] not driven (layer 3)
  // Warning: Z[53] not driven (layer 3)
  // Warning: Z[54] not driven (layer 3)
  // Warning: Z[55] not driven (layer 3)
  // Warning: Z[56] not driven (layer 3)
  // Warning: Z[57] not driven (layer 3)
  // Warning: Z[58] not driven (layer 3)
  // Warning: Z[59] not driven (layer 3)
  // Warning: Z[60] not driven (layer 3)
  // Warning: Z[61] not driven (layer 3)
  // Warning: Z[62] not driven (layer 3)
  // Warning: Z[63] not driven (layer 3)
  // Warning: Z[64] not driven (layer 3)
  // Warning: Z[65] not driven (layer 3)
  // Warning: Z[66] not driven (layer 3)
  // Warning: Z[67] not driven (layer 3)
  // Warning: Z[68] not driven (layer 3)
  // Warning: Z[69] not driven (layer 3)
  // Warning: Z[70] not driven (layer 3)
  // Warning: Z[71] not driven (layer 3)
  // Warning: Z[72] not driven (layer 3)
  // Warning: Z[73] not driven (layer 3)
  // Warning: Z[74] not driven (layer 3)
  // Warning: Z[75] not driven (layer 3)
  // Warning: Z[76] not driven (layer 3)
  // Warning: Z[77] not driven (layer 3)
  // Warning: Z[78] not driven (layer 3)
  // Warning: Z[79] not driven (layer 3)
  // Warning: Z[80] not driven (layer 3)
  // Warning: Z[81] not driven (layer 3)
  // Warning: Z[82] not driven (layer 3)
  // Warning: Z[83] not driven (layer 3)
  // Warning: Z[84] not driven (layer 3)
  // Warning: Z[85] not driven (layer 3)
  // Warning: Z[86] not driven (layer 3)
  // Warning: Z[87] not driven (layer 3)
  // Warning: Z[88] not driven (layer 3)
  // Warning: Z[89] not driven (layer 3)
  // Warning: Z[90] not driven (layer 3)
  // Warning: Z[91] not driven (layer 3)
  // Warning: Z[92] not driven (layer 3)
  // Warning: Z[93] not driven (layer 3)
  // Warning: Z[94] not driven (layer 3)
  // Warning: Z[95] not driven (layer 3)
  // Warning: Z[96] not driven (layer 3)
  // Warning: Z[97] not driven (layer 3)
  // Warning: Z[98] not driven (layer 3)
  // Warning: Z[99] not driven (layer 3)
  // Warning: Z[100] not driven (layer 3)
  // Warning: Z[101] not driven (layer 3)
  // Warning: Z[102] not driven (layer 3)
  // Warning: Z[103] not driven (layer 3)
  // Warning: Z[104] not driven (layer 3)
  // Warning: Z[105] not driven (layer 3)
  // Warning: Z[106] not driven (layer 3)
  // Warning: Z[107] not driven (layer 3)
  // Warning: Z[108] not driven (layer 3)
  // Warning: Z[109] not driven (layer 3)
  // Warning: Z[110] not driven (layer 3)
  // Warning: Z[111] not driven (layer 3)
  // Warning: Z[112] not driven (layer 3)
  // Warning: Z[113] not driven (layer 3)
  // Warning: Z[114] not driven (layer 3)
  // Warning: Z[115] not driven (layer 3)
  // Warning: Z[116] not driven (layer 3)
  // Warning: Z[117] not driven (layer 3)
  // Warning: Z[118] not driven (layer 3)
  // Warning: Z[119] not driven (layer 3)
  // Warning: Z[120] not driven (layer 3)
  // Warning: Z[121] not driven (layer 3)
  // Warning: Z[122] not driven (layer 3)
  // Warning: Z[123] not driven (layer 3)
  // Warning: Z[124] not driven (layer 3)
  // Warning: Z[125] not driven (layer 3)
  // Warning: Z[126] not driven (layer 3)
  // Warning: Z[127] not driven (layer 3)
  // Warning: Z[128] not driven (layer 3)
  // Warning: Z[129] not driven (layer 3)
  // Warning: Z[130] not driven (layer 3)
  // Warning: Z[131] not driven (layer 3)
  // Warning: Z[132] not driven (layer 3)
  // Warning: Z[133] not driven (layer 3)
  // Warning: Z[134] not driven (layer 3)
  // Warning: Z[135] not driven (layer 3)
  // Warning: Z[136] not driven (layer 3)
  // Warning: Z[137] not driven (layer 3)
  // Warning: Z[138] not driven (layer 3)
  // Warning: Z[139] not driven (layer 3)
  // Warning: Z[140] not driven (layer 3)
  // Warning: Z[141] not driven (layer 3)
  // Warning: Z[142] not driven (layer 3)
  // Warning: Z[143] not driven (layer 3)
  // Warning: Z[144] not driven (layer 3)
  // Warning: Z[145] not driven (layer 3)
  // Warning: Z[146] not driven (layer 3)
  // Warning: Z[147] not driven (layer 3)
  // Warning: Z[148] not driven (layer 3)
  // Warning: Z[149] not driven (layer 3)
  // Warning: Z[150] not driven (layer 3)
  // Warning: Z[151] not driven (layer 3)
  // Warning: Z[152] not driven (layer 3)
  // Warning: Z[153] not driven (layer 3)
  // Warning: Z[154] not driven (layer 3)
  // Warning: Z[155] not driven (layer 3)
  // Warning: Z[156] not driven (layer 3)
  // Warning: Z[157] not driven (layer 3)
  // Warning: Z[158] not driven (layer 3)
  // Warning: Z[159] not driven (layer 3)
  // Warning: Z[160] not driven (layer 3)
  // Warning: Z[161] not driven (layer 3)
  // Warning: Z[162] not driven (layer 3)
  // Warning: Z[163] not driven (layer 3)
  // Warning: Z[164] not driven (layer 3)
  // Warning: Z[165] not driven (layer 3)
  // Warning: Z[166] not driven (layer 3)
  // Warning: Z[167] not driven (layer 3)
  // Warning: Z[168] not driven (layer 3)
  // Warning: Z[169] not driven (layer 3)
  // Warning: Z[170] not driven (layer 3)
  // Warning: Z[171] not driven (layer 3)
  // Warning: Z[172] not driven (layer 3)
  // Warning: Z[173] not driven (layer 3)
  // Warning: Z[174] not driven (layer 3)
  // Warning: Z[175] not driven (layer 3)
  // Warning: Z[176] not driven (layer 3)
  // Warning: Z[177] not driven (layer 3)
  // Warning: Z[178] not driven (layer 3)
  // Warning: Z[179] not driven (layer 3)
  // Warning: Z[180] not driven (layer 3)
  // Warning: Z[181] not driven (layer 3)
  // Warning: Z[182] not driven (layer 3)
  // Warning: Z[183] not driven (layer 3)
  // Warning: Z[184] not driven (layer 3)
  // Warning: Z[185] not driven (layer 3)
  // Warning: Z[186] not driven (layer 3)
  // Warning: Z[187] not driven (layer 3)
  // Warning: Z[188] not driven (layer 3)
  // Warning: Z[189] not driven (layer 3)
  // Warning: Z[190] not driven (layer 3)
  // Warning: Z[191] not driven (layer 3)
  // Warning: Z[192] not driven (layer 3)
  // Warning: Z[193] not driven (layer 3)
  // Warning: Z[194] not driven (layer 3)
  // Warning: Z[195] not driven (layer 3)
  // Warning: Z[196] not driven (layer 3)
  // Warning: Z[197] not driven (layer 3)
  // Warning: Z[198] not driven (layer 3)
  // Warning: Z[199] not driven (layer 3)
  // Warning: Z[200] not driven (layer 3)
  // Warning: Z[201] not driven (layer 3)
  // Warning: Z[202] not driven (layer 3)
  // Warning: Z[203] not driven (layer 3)
  // Warning: Z[204] not driven (layer 3)
  // Warning: Z[205] not driven (layer 3)
  // Warning: Z[206] not driven (layer 3)
  // Warning: Z[207] not driven (layer 3)
  // Warning: Z[208] not driven (layer 3)
  // Warning: Z[209] not driven (layer 3)
  // Warning: Z[210] not driven (layer 3)
  // Warning: Z[211] not driven (layer 3)
  // Warning: Z[212] not driven (layer 3)
  // Warning: Z[213] not driven (layer 3)
  // Warning: Z[214] not driven (layer 3)
  // Warning: Z[215] not driven (layer 3)
  // Warning: Z[216] not driven (layer 3)
  // Warning: Z[217] not driven (layer 3)
  // Warning: Z[218] not driven (layer 3)
  // Warning: Z[219] not driven (layer 3)
  // Warning: Z[220] not driven (layer 3)
  // Warning: Z[221] not driven (layer 3)
  // Warning: Z[222] not driven (layer 3)
  // Warning: Z[223] not driven (layer 3)
  // Warning: Z[224] not driven (layer 3)
  // Warning: Z[225] not driven (layer 3)
  // Warning: Z[226] not driven (layer 3)
  // Warning: Z[227] not driven (layer 3)
  // Warning: Z[228] not driven (layer 3)
  // Warning: Z[229] not driven (layer 3)
  // Warning: Z[230] not driven (layer 3)
  // Warning: Z[231] not driven (layer 3)
  // Warning: Z[232] not driven (layer 3)
  // Warning: Z[233] not driven (layer 3)
  // Warning: Z[234] not driven (layer 3)
  // Warning: Z[235] not driven (layer 3)
  // Warning: Z[236] not driven (layer 3)
  // Warning: Z[237] not driven (layer 3)
  // Warning: Z[238] not driven (layer 3)
  // Warning: Z[239] not driven (layer 3)
  // Warning: Z[240] not driven (layer 3)
  // Warning: Z[241] not driven (layer 3)
  // Warning: Z[242] not driven (layer 3)
  // Warning: Z[243] not driven (layer 3)
  // Warning: Z[244] not driven (layer 3)
  // Warning: Z[245] not driven (layer 3)
  // Warning: Z[246] not driven (layer 3)
  // Warning: Z[247] not driven (layer 3)
  // Warning: Z[248] not driven (layer 3)
  // Warning: Z[249] not driven (layer 3)
  // Warning: Z[250] not driven (layer 3)
  // Warning: Z[251] not driven (layer 3)
  // Warning: Z[252] not driven (layer 3)
  // Warning: Z[253] not driven (layer 3)
  // Warning: Z[254] not driven (layer 3)
  // Warning: Z[255] not driven (layer 3)

endmodule
