`timescale 1ns / 1ps
`include "all_cmos_tf_rst_mnist.v"
`include "all_cmos_tf_rst.v"

module mnist_neural_network(
    input wire clk,
    input wire rst,
    input wire [115:0] input_layer, // TODO: widen if needed
    output wire [255:0] Z
);

  // Internal signals
  wire [255:0] Y; // layer 1 outputs feed layer 3

  // instantiate function_0 for neuron0_1
  function_0 neuron0_1 (
      .a(input_layer[541]),
      .b(input_layer[1947]),
      .c(input_layer[1804]),
      .d(~input_layer[537]),
      .e(~input_layer[1985]),
      .y(Y[0]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1_1
  function_1 neuron1_1 (
      .a(~input_layer[715]),
      .b(~input_layer[2220]),
      .c(~input_layer[1790]),
      .d(~input_layer[371]),
      .e(~input_layer[1634]),
      .f(input_layer[2138]),
      .y(Y[1]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_2 for neuron2_1
  function_2 neuron2_1 (
      .a(input_layer[1272]),
      .b(input_layer[739]),
      .c(~input_layer[1066]),
      .d(input_layer[1417]),
      .e(input_layer[1652]),
      .f(input_layer[71]),
      .y(Y[2]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron3_1
  function_3 neuron3_1 (
      .a(input_layer[2133]),
      .b(input_layer[497]),
      .c(input_layer[1276]),
      .d(~input_layer[553]),
      .e(input_layer[482]),
      .y(Y[3]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron4_1
  function_4 neuron4_1 (
      .a(input_layer[1973]),
      .b(~input_layer[379]),
      .c(input_layer[1967]),
      .d(~input_layer[1607]),
      .e(~input_layer[1556]),
      .y(Y[4]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron5_1
  function_5 neuron5_1 (
      .a(input_layer[819]),
      .b(input_layer[2131]),
      .y(Y[5]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron6_1
  function_6 neuron6_1 (
      .a(~input_layer[964]),
      .b(input_layer[1610]),
      .c(input_layer[1214]),
      .d(~input_layer[1574]),
      .e(input_layer[1177]),
      .f(input_layer[1516]),
      .y(Y[6]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron7_1
  function_7 neuron7_1 (
      .a(input_layer[463]),
      .b(~input_layer[125]),
      .c(input_layer[1835]),
      .d(input_layer[1648]),
      .e(input_layer[1856]),
      .f(input_layer[1031]),
      .y(Y[7]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron8_1
  function_8 neuron8_1 (
      .a(~input_layer[1832]),
      .b(~input_layer[523]),
      .c(~input_layer[639]),
      .d(input_layer[926]),
      .e(input_layer[1599]),
      .f(input_layer[1431]),
      .y(Y[8]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_9 for neuron9_1
  function_9 neuron9_1 (
      .a(~input_layer[1134]),
      .b(input_layer[1539]),
      .c(~input_layer[467]),
      .d(~input_layer[2232]),
      .e(input_layer[866]),
      .y(Y[9]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron10_1
  function_10 neuron10_1 (
      .a(~input_layer[1216]),
      .b(input_layer[137]),
      .c(~input_layer[946]),
      .d(input_layer[367]),
      .y(Y[10]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron11_1
  function_11 neuron11_1 (
      .a(input_layer[2236]),
      .b(input_layer[2144]),
      .c(input_layer[1626]),
      .d(input_layer[1859]),
      .y(Y[11]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron12_1
  function_12 neuron12_1 (
      .a(~input_layer[1143]),
      .b(~input_layer[778]),
      .c(~input_layer[639]),
      .y(Y[12]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron13_1
  function_13 neuron13_1 (
      .a(~input_layer[1701]),
      .b(input_layer[1154]),
      .c(~input_layer[1730]),
      .d(input_layer[2074]),
      .e(input_layer[1964]),
      .f(input_layer[2214]),
      .y(Y[13]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron14_1
  function_14 neuron14_1 (
      .a(~input_layer[1208]),
      .b(~input_layer[2209]),
      .c(~input_layer[670]),
      .d(input_layer[2008]),
      .e(~input_layer[155]),
      .y(Y[14]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_15 for neuron15_1
  function_15 neuron15_1 (
      .a(~input_layer[1378]),
      .b(~input_layer[1631]),
      .c(input_layer[1167]),
      .d(~input_layer[1223]),
      .e(input_layer[978]),
      .f(input_layer[1107]),
      .y(Y[15]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron16_1
  function_16 neuron16_1 (
      .a(input_layer[830]),
      .b(input_layer[354]),
      .c(input_layer[597]),
      .y(Y[16]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[17] = 1'b0;

  // instantiate function_17 for neuron18_1
  function_17 neuron18_1 (
      .a(~input_layer[1780]),
      .b(~input_layer[1785]),
      .c(input_layer[1484]),
      .d(~input_layer[764]),
      .e(~input_layer[2201]),
      .f(~input_layer[2004]),
      .y(Y[18]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron19_1
  function_18 neuron19_1 (
      .a(~input_layer[1354]),
      .b(input_layer[1706]),
      .c(~input_layer[1236]),
      .d(~input_layer[2327]),
      .e(~input_layer[1647]),
      .y(Y[19]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron20_1
  function_19 neuron20_1 (
      .a(~input_layer[449]),
      .b(input_layer[1123]),
      .c(~input_layer[1216]),
      .d(input_layer[2290]),
      .y(Y[20]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron21_1
  function_20 neuron21_1 (
      .a(input_layer[1160]),
      .b(input_layer[1979]),
      .c(input_layer[738]),
      .d(~input_layer[1152]),
      .e(input_layer[1274]),
      .f(~input_layer[1374]),
      .y(Y[21]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron22_1
  function_21 neuron22_1 (
      .a(~input_layer[1561]),
      .b(~input_layer[959]),
      .c(~input_layer[520]),
      .d(~input_layer[2174]),
      .y(Y[22]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron23_1
  function_18 neuron23_1 (
      .a(~input_layer[1446]),
      .b(~input_layer[395]),
      .c(~input_layer[312]),
      .d(~input_layer[196]),
      .e(~input_layer[1443]),
      .y(Y[23]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron24_1
  function_18 neuron24_1 (
      .a(~input_layer[1032]),
      .b(input_layer[785]),
      .c(~input_layer[2026]),
      .d(~input_layer[443]),
      .e(~input_layer[2088]),
      .y(Y[24]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_22 for neuron25_1
  function_22 neuron25_1 (
      .a(~input_layer[1611]),
      .b(input_layer[486]),
      .c(~input_layer[694]),
      .d(~input_layer[512]),
      .e(input_layer[1433]),
      .f(~input_layer[1684]),
      .y(Y[25]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_23 for neuron26_1
  function_23 neuron26_1 (
      .a(input_layer[846]),
      .b(~input_layer[1384]),
      .c(~input_layer[1296]),
      .d(~input_layer[595]),
      .e(~input_layer[2108]),
      .f(~input_layer[1910]),
      .y(Y[26]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron27_1
  function_24 neuron27_1 (
      .a(input_layer[1188]),
      .y(Y[27]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron28_1
  function_16 neuron28_1 (
      .a(input_layer[1854]),
      .b(input_layer[655]),
      .c(input_layer[637]),
      .y(Y[28]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron29_1
  function_25 neuron29_1 (
      .a(input_layer[403]),
      .b(input_layer[2080]),
      .c(input_layer[2202]),
      .d(input_layer[2320]),
      .e(~input_layer[1293]),
      .y(Y[29]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron30_1
  function_26 neuron30_1 (
      .a(~input_layer[1231]),
      .b(~input_layer[1806]),
      .y(Y[30]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_27 for neuron31_1
  function_27 neuron31_1 (
      .a(input_layer[1165]),
      .b(~input_layer[1104]),
      .c(input_layer[1665]),
      .d(input_layer[1739]),
      .e(~input_layer[2073]),
      .f(input_layer[456]),
      .y(Y[31]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron32_1
  function_28 neuron32_1 (
      .a(input_layer[573]),
      .b(input_layer[823]),
      .c(~input_layer[283]),
      .d(~input_layer[537]),
      .e(input_layer[677]),
      .f(~input_layer[1342]),
      .y(Y[32]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron33_1
  function_29 neuron33_1 (
      .a(~input_layer[489]),
      .b(input_layer[1360]),
      .c(input_layer[1276]),
      .d(~input_layer[1986]),
      .e(~input_layer[1766]),
      .f(input_layer[13]),
      .y(Y[33]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron34_1
  function_30 neuron34_1 (
      .a(input_layer[1774]),
      .b(~input_layer[1196]),
      .c(input_layer[430]),
      .d(~input_layer[1105]),
      .y(Y[34]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron35_1
  function_21 neuron35_1 (
      .a(~input_layer[298]),
      .b(~input_layer[436]),
      .c(~input_layer[1078]),
      .d(~input_layer[109]),
      .y(Y[35]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron36_1
  function_31 neuron36_1 (
      .a(input_layer[1746]),
      .b(input_layer[137]),
      .c(input_layer[111]),
      .d(input_layer[2010]),
      .e(~input_layer[539]),
      .f(input_layer[2280]),
      .y(Y[36]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron37_1
  function_14 neuron37_1 (
      .a(~input_layer[232]),
      .b(input_layer[664]),
      .c(~input_layer[2299]),
      .d(input_layer[656]),
      .e(input_layer[1988]),
      .y(Y[37]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron38_1
  function_32 neuron38_1 (
      .a(~input_layer[1813]),
      .b(input_layer[2035]),
      .c(input_layer[1675]),
      .d(input_layer[1927]),
      .y(Y[38]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron39_1
  function_33 neuron39_1 (
      .a(~input_layer[2203]),
      .b(~input_layer[682]),
      .c(~input_layer[958]),
      .d(~input_layer[1288]),
      .e(input_layer[183]),
      .y(Y[39]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron40_1
  function_34 neuron40_1 (
      .a(~input_layer[1053]),
      .b(input_layer[302]),
      .c(input_layer[1631]),
      .d(input_layer[1623]),
      .e(input_layer[1414]),
      .y(Y[40]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron41_1
  function_33 neuron41_1 (
      .a(~input_layer[223]),
      .b(~input_layer[1915]),
      .c(~input_layer[203]),
      .d(~input_layer[1116]),
      .e(input_layer[1939]),
      .y(Y[41]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron42_1
  function_0 neuron42_1 (
      .a(input_layer[851]),
      .b(input_layer[271]),
      .c(input_layer[460]),
      .d(input_layer[2035]),
      .e(~input_layer[949]),
      .y(Y[42]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron43_1
  function_35 neuron43_1 (
      .a(~input_layer[604]),
      .b(input_layer[315]),
      .c(~input_layer[550]),
      .d(~input_layer[355]),
      .e(~input_layer[2111]),
      .y(Y[43]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron44_1
  function_36 neuron44_1 (
      .a(input_layer[918]),
      .b(~input_layer[1240]),
      .c(~input_layer[930]),
      .d(input_layer[1949]),
      .e(input_layer[777]),
      .f(input_layer[779]),
      .y(Y[44]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron45_1
  function_0 neuron45_1 (
      .a(input_layer[1295]),
      .b(input_layer[1376]),
      .c(input_layer[1139]),
      .d(input_layer[1507]),
      .e(input_layer[1045]),
      .y(Y[45]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron46_1
  function_37 neuron46_1 (
      .a(input_layer[1557]),
      .b(~input_layer[2141]),
      .c(input_layer[1273]),
      .d(~input_layer[463]),
      .e(input_layer[1081]),
      .y(Y[46]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron47_1
  function_16 neuron47_1 (
      .a(input_layer[463]),
      .b(input_layer[1335]),
      .c(input_layer[1923]),
      .y(Y[47]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron48_1
  function_3 neuron48_1 (
      .a(input_layer[1280]),
      .b(input_layer[1607]),
      .c(input_layer[2124]),
      .d(~input_layer[419]),
      .e(~input_layer[990]),
      .y(Y[48]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_38 for neuron49_1
  function_38 neuron49_1 (
      .a(input_layer[1457]),
      .b(~input_layer[1864]),
      .c(input_layer[399]),
      .d(input_layer[1173]),
      .e(input_layer[2177]),
      .f(input_layer[1229]),
      .y(Y[49]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron50_1
  function_39 neuron50_1 (
      .a(input_layer[531]),
      .b(~input_layer[576]),
      .c(~input_layer[1878]),
      .d(input_layer[1617]),
      .y(Y[50]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron51_1
  function_40 neuron51_1 (
      .a(~input_layer[606]),
      .b(~input_layer[1855]),
      .c(input_layer[1791]),
      .d(~input_layer[429]),
      .e(input_layer[1071]),
      .f(~input_layer[1013]),
      .y(Y[51]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_41 for neuron52_1
  function_41 neuron52_1 (
      .a(input_layer[447]),
      .b(input_layer[1329]),
      .c(~input_layer[1185]),
      .d(~input_layer[2220]),
      .e(input_layer[1537]),
      .f(~input_layer[2198]),
      .y(Y[52]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron53_1
  function_3 neuron53_1 (
      .a(input_layer[1127]),
      .b(input_layer[1611]),
      .c(input_layer[438]),
      .d(~input_layer[978]),
      .e(input_layer[1148]),
      .y(Y[53]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron54_1
  function_42 neuron54_1 (
      .a(~input_layer[1551]),
      .b(input_layer[395]),
      .c(~input_layer[1461]),
      .d(~input_layer[417]),
      .e(~input_layer[1852]),
      .y(Y[54]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron55_1
  function_43 neuron55_1 (
      .a(input_layer[1423]),
      .b(~input_layer[500]),
      .c(~input_layer[1133]),
      .d(input_layer[439]),
      .e(~input_layer[679]),
      .y(Y[55]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron56_1
  function_44 neuron56_1 (
      .a(~input_layer[1138]),
      .b(~input_layer[2051]),
      .c(~input_layer[916]),
      .y(Y[56]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron57_1
  function_14 neuron57_1 (
      .a(~input_layer[2203]),
      .b(input_layer[1881]),
      .c(~input_layer[2164]),
      .d(~input_layer[121]),
      .e(~input_layer[1003]),
      .y(Y[57]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron58_1
  function_34 neuron58_1 (
      .a(input_layer[1821]),
      .b(input_layer[1522]),
      .c(~input_layer[1231]),
      .d(~input_layer[1404]),
      .e(input_layer[1359]),
      .y(Y[58]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron59_1
  function_45 neuron59_1 (
      .a(~input_layer[1325]),
      .b(~input_layer[2202]),
      .c(~input_layer[239]),
      .d(~input_layer[1058]),
      .e(~input_layer[471]),
      .f(~input_layer[1180]),
      .y(Y[59]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_46 for neuron60_1
  function_46 neuron60_1 (
      .a(input_layer[2228]),
      .b(~input_layer[1300]),
      .c(~input_layer[1422]),
      .d(input_layer[356]),
      .e(input_layer[1194]),
      .f(input_layer[104]),
      .y(Y[60]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron61_1
  function_5 neuron61_1 (
      .a(~input_layer[1204]),
      .b(input_layer[1005]),
      .y(Y[61]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron62_1
  function_18 neuron62_1 (
      .a(~input_layer[2174]),
      .b(input_layer[368]),
      .c(input_layer[373]),
      .d(~input_layer[1208]),
      .e(~input_layer[2041]),
      .y(Y[62]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron63_1
  function_26 neuron63_1 (
      .a(~input_layer[225]),
      .b(~input_layer[946]),
      .y(Y[63]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_47 for neuron64_1
  function_47 neuron64_1 (
      .a(~input_layer[1130]),
      .b(~input_layer[1367]),
      .c(input_layer[2168]),
      .d(~input_layer[201]),
      .e(~input_layer[361]),
      .f(input_layer[1541]),
      .y(Y[64]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron65_1
  function_48 neuron65_1 (
      .a(input_layer[2323]),
      .b(~input_layer[982]),
      .c(~input_layer[2223]),
      .d(input_layer[2217]),
      .e(input_layer[1257]),
      .y(Y[65]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron66_1
  function_49 neuron66_1 (
      .a(input_layer[1161]),
      .b(input_layer[121]),
      .c(input_layer[690]),
      .d(input_layer[774]),
      .e(input_layer[2173]),
      .f(input_layer[1492]),
      .y(Y[66]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_50 for neuron67_1
  function_50 neuron67_1 (
      .a(~input_layer[2138]),
      .b(~input_layer[1745]),
      .c(input_layer[1418]),
      .d(~input_layer[1089]),
      .e(input_layer[150]),
      .y(Y[67]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_51 for neuron68_1
  function_51 neuron68_1 (
      .a(input_layer[2046]),
      .b(input_layer[1840]),
      .c(input_layer[681]),
      .d(~input_layer[1334]),
      .e(input_layer[1172]),
      .f(~input_layer[867]),
      .y(Y[68]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron69_1
  function_52 neuron69_1 (
      .a(~input_layer[141]),
      .b(input_layer[1155]),
      .c(~input_layer[2052]),
      .d(~input_layer[1883]),
      .e(input_layer[323]),
      .y(Y[69]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron70_1
  function_16 neuron70_1 (
      .a(input_layer[947]),
      .b(input_layer[912]),
      .c(~input_layer[365]),
      .y(Y[70]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron71_1
  function_53 neuron71_1 (
      .a(input_layer[2159]),
      .b(~input_layer[693]),
      .c(input_layer[1440]),
      .d(input_layer[2012]),
      .e(input_layer[74]),
      .y(Y[71]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron72_1
  function_35 neuron72_1 (
      .a(~input_layer[524]),
      .b(~input_layer[1076]),
      .c(input_layer[738]),
      .d(~input_layer[1359]),
      .e(~input_layer[1456]),
      .y(Y[72]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron73_1
  function_10 neuron73_1 (
      .a(input_layer[818]),
      .b(input_layer[1021]),
      .c(~input_layer[316]),
      .d(input_layer[2201]),
      .y(Y[73]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron74_1
  function_54 neuron74_1 (
      .a(input_layer[2241]),
      .b(input_layer[228]),
      .c(input_layer[1171]),
      .d(~input_layer[1324]),
      .e(~input_layer[690]),
      .f(input_layer[1565]),
      .y(Y[74]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron75_1
  function_55 neuron75_1 (
      .a(input_layer[1407]),
      .b(~input_layer[141]),
      .c(~input_layer[1128]),
      .d(~input_layer[1243]),
      .e(input_layer[1071]),
      .f(input_layer[1621]),
      .y(Y[75]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron76_1
  function_56 neuron76_1 (
      .a(~input_layer[1714]),
      .b(~input_layer[116]),
      .c(~input_layer[307]),
      .d(input_layer[1203]),
      .e(~input_layer[1648]),
      .y(Y[76]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_57 for neuron77_1
  function_57 neuron77_1 (
      .a(~input_layer[2311]),
      .b(input_layer[489]),
      .c(~input_layer[900]),
      .d(input_layer[1476]),
      .e(~input_layer[453]),
      .f(input_layer[1209]),
      .y(Y[77]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_58 for neuron78_1
  function_58 neuron78_1 (
      .a(~input_layer[824]),
      .b(~input_layer[690]),
      .c(input_layer[147]),
      .d(input_layer[1157]),
      .e(input_layer[990]),
      .f(~input_layer[355]),
      .y(Y[78]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron79_1
  function_32 neuron79_1 (
      .a(input_layer[1580]),
      .b(input_layer[454]),
      .c(~input_layer[597]),
      .d(input_layer[1367]),
      .y(Y[79]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron80_1
  function_11 neuron80_1 (
      .a(input_layer[1722]),
      .b(input_layer[204]),
      .c(input_layer[1602]),
      .d(~input_layer[702]),
      .y(Y[80]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron81_1
  function_16 neuron81_1 (
      .a(input_layer[610]),
      .b(input_layer[1773]),
      .c(input_layer[1442]),
      .y(Y[81]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron82_1
  function_25 neuron82_1 (
      .a(input_layer[915]),
      .b(input_layer[325]),
      .c(input_layer[745]),
      .d(input_layer[1411]),
      .e(input_layer[683]),
      .y(Y[82]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron83_1
  function_59 neuron83_1 (
      .a(~input_layer[1585]),
      .b(~input_layer[1716]),
      .c(~input_layer[604]),
      .d(input_layer[1311]),
      .e(input_layer[1353]),
      .f(input_layer[1999]),
      .y(Y[83]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron84_1
  function_60 neuron84_1 (
      .a(~input_layer[329]),
      .b(input_layer[1707]),
      .c(~input_layer[777]),
      .d(~input_layer[131]),
      .e(input_layer[903]),
      .f(~input_layer[300]),
      .y(Y[84]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron85_1
  function_14 neuron85_1 (
      .a(~input_layer[1250]),
      .b(input_layer[1216]),
      .c(~input_layer[1427]),
      .d(~input_layer[1741]),
      .e(~input_layer[1883]),
      .y(Y[85]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron86_1
  function_35 neuron86_1 (
      .a(~input_layer[1288]),
      .b(~input_layer[1504]),
      .c(~input_layer[1079]),
      .d(input_layer[1102]),
      .e(input_layer[426]),
      .y(Y[86]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron87_1
  function_61 neuron87_1 (
      .a(~input_layer[438]),
      .b(~input_layer[533]),
      .c(~input_layer[2177]),
      .d(~input_layer[1429]),
      .e(input_layer[2071]),
      .y(Y[87]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron88_1
  function_48 neuron88_1 (
      .a(input_layer[1835]),
      .b(~input_layer[529]),
      .c(input_layer[1011]),
      .d(~input_layer[1136]),
      .e(~input_layer[1567]),
      .y(Y[88]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron89_1
  function_62 neuron89_1 (
      .a(~input_layer[1478]),
      .b(~input_layer[1440]),
      .c(input_layer[1872]),
      .d(~input_layer[1994]),
      .y(Y[89]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron90_1
  function_34 neuron90_1 (
      .a(input_layer[2050]),
      .b(input_layer[763]),
      .c(input_layer[512]),
      .d(~input_layer[1398]),
      .e(~input_layer[1844]),
      .y(Y[90]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron91_1
  function_63 neuron91_1 (
      .a(input_layer[1925]),
      .b(~input_layer[1989]),
      .c(~input_layer[471]),
      .d(~input_layer[1054]),
      .y(Y[91]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron92_1
  function_1 neuron92_1 (
      .a(~input_layer[1451]),
      .b(~input_layer[2147]),
      .c(~input_layer[927]),
      .d(input_layer[1704]),
      .e(~input_layer[1655]),
      .f(input_layer[966]),
      .y(Y[92]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron93_1
  function_64 neuron93_1 (
      .a(input_layer[831]),
      .b(input_layer[288]),
      .c(~input_layer[1289]),
      .d(input_layer[1481]),
      .e(~input_layer[700]),
      .y(Y[93]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron94_1
  function_11 neuron94_1 (
      .a(input_layer[2152]),
      .b(input_layer[2220]),
      .c(input_layer[1944]),
      .d(~input_layer[1458]),
      .y(Y[94]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron95_1
  function_26 neuron95_1 (
      .a(input_layer[2320]),
      .b(~input_layer[1605]),
      .y(Y[95]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron96_1
  function_65 neuron96_1 (
      .a(~input_layer[1876]),
      .b(~input_layer[2315]),
      .c(input_layer[1158]),
      .d(input_layer[203]),
      .e(input_layer[1140]),
      .f(~input_layer[1897]),
      .y(Y[96]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_66 for neuron97_1
  function_66 neuron97_1 (
      .a(~input_layer[455]),
      .b(input_layer[2301]),
      .c(~input_layer[620]),
      .d(~input_layer[1962]),
      .e(~input_layer[2325]),
      .f(input_layer[107]),
      .y(Y[97]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron98_1
  function_67 neuron98_1 (
      .a(input_layer[1783]),
      .b(input_layer[1015]),
      .c(~input_layer[1201]),
      .d(~input_layer[2084]),
      .e(input_layer[1805]),
      .y(Y[98]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron99_1
  function_43 neuron99_1 (
      .a(input_layer[797]),
      .b(~input_layer[1909]),
      .c(~input_layer[1823]),
      .d(~input_layer[1559]),
      .e(~input_layer[535]),
      .y(Y[99]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_68 for neuron100_1
  function_68 neuron100_1 (
      .a(~input_layer[912]),
      .b(input_layer[1775]),
      .c(~input_layer[1540]),
      .d(~input_layer[823]),
      .e(~input_layer[1211]),
      .f(input_layer[74]),
      .y(Y[100]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron101_1
  function_11 neuron101_1 (
      .a(input_layer[1585]),
      .b(input_layer[374]),
      .c(input_layer[1520]),
      .d(input_layer[700]),
      .y(Y[101]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron102_1
  function_69 neuron102_1 (
      .a(input_layer[799]),
      .b(input_layer[2125]),
      .c(~input_layer[1806]),
      .d(~input_layer[962]),
      .e(input_layer[1260]),
      .y(Y[102]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron103_1
  function_70 neuron103_1 (
      .a(~input_layer[894]),
      .b(input_layer[1536]),
      .c(~input_layer[2253]),
      .d(input_layer[265]),
      .e(input_layer[63]),
      .f(input_layer[2020]),
      .y(Y[103]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron104_1
  function_37 neuron104_1 (
      .a(~input_layer[717]),
      .b(input_layer[1990]),
      .c(input_layer[306]),
      .d(~input_layer[2140]),
      .e(~input_layer[784]),
      .y(Y[104]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_71 for neuron105_1
  function_71 neuron105_1 (
      .a(input_layer[1326]),
      .b(input_layer[220]),
      .c(input_layer[1239]),
      .d(~input_layer[1095]),
      .e(~input_layer[1096]),
      .f(~input_layer[1174]),
      .y(Y[105]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron106_1
  function_25 neuron106_1 (
      .a(input_layer[613]),
      .b(input_layer[542]),
      .c(input_layer[773]),
      .d(input_layer[1604]),
      .e(input_layer[1943]),
      .y(Y[106]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron107_1
  function_72 neuron107_1 (
      .a(~input_layer[1156]),
      .b(~input_layer[1317]),
      .c(input_layer[2216]),
      .d(~input_layer[2131]),
      .e(input_layer[1593]),
      .y(Y[107]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_73 for neuron108_1
  function_73 neuron108_1 (
      .a(input_layer[2135]),
      .b(~input_layer[1903]),
      .c(~input_layer[1961]),
      .d(input_layer[1732]),
      .e(~input_layer[2070]),
      .f(input_layer[99]),
      .y(Y[108]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron109_1
  function_74 neuron109_1 (
      .a(input_layer[2126]),
      .b(~input_layer[349]),
      .c(~input_layer[1876]),
      .d(input_layer[687]),
      .e(~input_layer[1073]),
      .y(Y[109]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron110_1
  function_75 neuron110_1 (
      .a(~input_layer[1668]),
      .b(~input_layer[1917]),
      .c(input_layer[209]),
      .d(input_layer[1686]),
      .e(~input_layer[1250]),
      .y(Y[110]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron111_1
  function_5 neuron111_1 (
      .a(input_layer[311]),
      .b(~input_layer[1629]),
      .y(Y[111]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron112_1
  function_11 neuron112_1 (
      .a(input_layer[391]),
      .b(input_layer[1414]),
      .c(input_layer[684]),
      .d(input_layer[1874]),
      .y(Y[112]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron113_1
  function_76 neuron113_1 (
      .a(~input_layer[1458]),
      .b(~input_layer[742]),
      .c(~input_layer[659]),
      .d(~input_layer[122]),
      .e(input_layer[1192]),
      .f(input_layer[1239]),
      .y(Y[113]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron114_1
  function_35 neuron114_1 (
      .a(~input_layer[819]),
      .b(~input_layer[813]),
      .c(~input_layer[1840]),
      .d(~input_layer[457]),
      .e(input_layer[426]),
      .y(Y[114]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_77 for neuron115_1
  function_77 neuron115_1 (
      .a(~input_layer[217]),
      .b(input_layer[943]),
      .c(input_layer[1975]),
      .d(input_layer[837]),
      .e(input_layer[1312]),
      .f(input_layer[982]),
      .y(Y[115]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_78 for neuron116_1
  function_78 neuron116_1 (
      .a(input_layer[1468]),
      .b(input_layer[1854]),
      .c(~input_layer[1446]),
      .d(~input_layer[1166]),
      .e(input_layer[1691]),
      .f(~input_layer[1492]),
      .y(Y[116]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_79 for neuron117_1
  function_79 neuron117_1 (
      .a(~input_layer[1530]),
      .b(~input_layer[1819]),
      .c(input_layer[1942]),
      .d(input_layer[1808]),
      .e(~input_layer[1564]),
      .f(~input_layer[1709]),
      .y(Y[117]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_80 for neuron118_1
  function_80 neuron118_1 (
      .a(~input_layer[1204]),
      .b(input_layer[1897]),
      .c(~input_layer[1394]),
      .d(input_layer[1979]),
      .e(input_layer[523]),
      .f(input_layer[1020]),
      .y(Y[118]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron119_1
  function_67 neuron119_1 (
      .a(input_layer[289]),
      .b(input_layer[2121]),
      .c(~input_layer[2060]),
      .d(input_layer[1516]),
      .e(~input_layer[612]),
      .y(Y[119]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron120_1
  function_35 neuron120_1 (
      .a(~input_layer[2322]),
      .b(input_layer[1285]),
      .c(~input_layer[2217]),
      .d(input_layer[2240]),
      .e(~input_layer[1087]),
      .y(Y[120]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_81 for neuron121_1
  function_81 neuron121_1 (
      .a(~input_layer[1362]),
      .b(input_layer[885]),
      .c(~input_layer[2050]),
      .d(input_layer[2094]),
      .e(input_layer[1697]),
      .f(~input_layer[1929]),
      .y(Y[121]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron122_1
  function_26 neuron122_1 (
      .a(~input_layer[1686]),
      .b(~input_layer[456]),
      .y(Y[122]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron123_1
  function_72 neuron123_1 (
      .a(~input_layer[1053]),
      .b(input_layer[1047]),
      .c(~input_layer[1272]),
      .d(input_layer[926]),
      .e(input_layer[716]),
      .y(Y[123]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron124_1
  function_82 neuron124_1 (
      .a(~input_layer[1700]),
      .b(input_layer[1064]),
      .c(input_layer[1357]),
      .d(~input_layer[1695]),
      .e(~input_layer[673]),
      .y(Y[124]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron125_1
  function_37 neuron125_1 (
      .a(input_layer[2316]),
      .b(~input_layer[1732]),
      .c(input_layer[671]),
      .d(input_layer[1378]),
      .e(~input_layer[1246]),
      .y(Y[125]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron126_1
  function_24 neuron126_1 (
      .a(input_layer[788]),
      .y(Y[126]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_83 for neuron127_1
  function_83 neuron127_1 (
      .a(input_layer[305]),
      .b(input_layer[1695]),
      .c(~input_layer[1049]),
      .d(~input_layer[1862]),
      .e(input_layer[1125]),
      .f(~input_layer[879]),
      .y(Y[127]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron128_1
  function_14 neuron128_1 (
      .a(~input_layer[1917]),
      .b(~input_layer[1420]),
      .c(~input_layer[502]),
      .d(~input_layer[670]),
      .e(~input_layer[669]),
      .y(Y[128]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron129_1
  function_24 neuron129_1 (
      .a(~input_layer[1221]),
      .y(Y[129]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron130_1
  function_84 neuron130_1 (
      .a(~input_layer[2231]),
      .b(~input_layer[2298]),
      .c(input_layer[1530]),
      .d(~input_layer[2332]),
      .e(input_layer[1734]),
      .f(input_layer[498]),
      .y(Y[130]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron131_1
  function_85 neuron131_1 (
      .a(input_layer[1548]),
      .b(input_layer[519]),
      .c(input_layer[2245]),
      .d(~input_layer[1539]),
      .e(~input_layer[1535]),
      .f(input_layer[2252]),
      .y(Y[131]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron132_1
  function_14 neuron132_1 (
      .a(~input_layer[1141]),
      .b(~input_layer[2003]),
      .c(~input_layer[1854]),
      .d(~input_layer[2012]),
      .e(~input_layer[1990]),
      .y(Y[132]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_86 for neuron133_1
  function_86 neuron133_1 (
      .a(input_layer[1528]),
      .b(input_layer[1961]),
      .c(input_layer[643]),
      .d(~input_layer[1604]),
      .e(~input_layer[118]),
      .f(~input_layer[988]),
      .y(Y[133]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron134_1
  function_18 neuron134_1 (
      .a(~input_layer[907]),
      .b(~input_layer[1393]),
      .c(~input_layer[769]),
      .d(~input_layer[2231]),
      .e(~input_layer[2205]),
      .y(Y[134]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_13 for neuron135_1
  function_13 neuron135_1 (
      .a(input_layer[1366]),
      .b(~input_layer[319]),
      .c(~input_layer[297]),
      .d(input_layer[2239]),
      .e(input_layer[569]),
      .f(~input_layer[1736]),
      .y(Y[135]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron136_1
  function_63 neuron136_1 (
      .a(input_layer[1861]),
      .b(~input_layer[1461]),
      .c(input_layer[272]),
      .d(~input_layer[1252]),
      .y(Y[136]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron137_1
  function_76 neuron137_1 (
      .a(~input_layer[446]),
      .b(~input_layer[1870]),
      .c(~input_layer[1222]),
      .d(~input_layer[121]),
      .e(~input_layer[1609]),
      .f(~input_layer[1733]),
      .y(Y[137]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron138_1
  function_43 neuron138_1 (
      .a(input_layer[1275]),
      .b(~input_layer[904]),
      .c(~input_layer[241]),
      .d(~input_layer[1969]),
      .e(~input_layer[176]),
      .y(Y[138]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron139_1
  function_12 neuron139_1 (
      .a(~input_layer[1732]),
      .b(~input_layer[1477]),
      .c(~input_layer[2084]),
      .y(Y[139]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron140_1
  function_87 neuron140_1 (
      .a(input_layer[1187]),
      .b(input_layer[1050]),
      .c(input_layer[268]),
      .d(input_layer[431]),
      .e(~input_layer[824]),
      .f(~input_layer[1875]),
      .y(Y[140]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron141_1
  function_40 neuron141_1 (
      .a(~input_layer[1972]),
      .b(~input_layer[196]),
      .c(~input_layer[752]),
      .d(~input_layer[210]),
      .e(~input_layer[409]),
      .f(~input_layer[1295]),
      .y(Y[141]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_88 for neuron142_1
  function_88 neuron142_1 (
      .a(input_layer[906]),
      .b(~input_layer[932]),
      .c(~input_layer[1255]),
      .d(~input_layer[1831]),
      .e(~input_layer[1736]),
      .f(~input_layer[753]),
      .y(Y[142]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron143_1
  function_89 neuron143_1 (
      .a(input_layer[1306]),
      .b(~input_layer[1451]),
      .c(~input_layer[1161]),
      .d(input_layer[2131]),
      .e(input_layer[1066]),
      .f(input_layer[1900]),
      .y(Y[143]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron144_1
  function_25 neuron144_1 (
      .a(input_layer[1062]),
      .b(input_layer[998]),
      .c(input_layer[314]),
      .d(input_layer[767]),
      .e(input_layer[416]),
      .y(Y[144]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron145_1
  function_90 neuron145_1 (
      .a(~input_layer[1165]),
      .b(~input_layer[1150]),
      .c(~input_layer[180]),
      .d(input_layer[812]),
      .e(~input_layer[1307]),
      .y(Y[145]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron146_1
  function_8 neuron146_1 (
      .a(~input_layer[1163]),
      .b(~input_layer[1025]),
      .c(input_layer[1738]),
      .d(input_layer[1588]),
      .e(~input_layer[808]),
      .f(input_layer[671]),
      .y(Y[146]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron147_1
  function_3 neuron147_1 (
      .a(input_layer[1812]),
      .b(input_layer[1455]),
      .c(~input_layer[706]),
      .d(input_layer[1561]),
      .e(input_layer[1007]),
      .y(Y[147]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron148_1
  function_21 neuron148_1 (
      .a(~input_layer[1590]),
      .b(~input_layer[107]),
      .c(input_layer[1808]),
      .d(~input_layer[2113]),
      .y(Y[148]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron149_1
  function_26 neuron149_1 (
      .a(input_layer[957]),
      .b(input_layer[564]),
      .y(Y[149]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron150_1
  function_24 neuron150_1 (
      .a(~input_layer[1283]),
      .y(Y[150]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[151] = 1'b0;

  // instantiate function_91 for neuron152_1
  function_91 neuron152_1 (
      .a(input_layer[1078]),
      .b(input_layer[1064]),
      .c(~input_layer[655]),
      .d(input_layer[1351]),
      .e(input_layer[174]),
      .f(~input_layer[949]),
      .y(Y[152]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron153_1
  function_92 neuron153_1 (
      .a(~input_layer[833]),
      .b(input_layer[977]),
      .c(input_layer[1357]),
      .d(~input_layer[410]),
      .y(Y[153]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron154_1
  function_16 neuron154_1 (
      .a(input_layer[1964]),
      .b(input_layer[1796]),
      .c(input_layer[624]),
      .y(Y[154]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron155_1
  function_3 neuron155_1 (
      .a(input_layer[229]),
      .b(input_layer[317]),
      .c(input_layer[1940]),
      .d(~input_layer[1797]),
      .e(~input_layer[1495]),
      .y(Y[155]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron156_1
  function_93 neuron156_1 (
      .a(~input_layer[997]),
      .b(~input_layer[766]),
      .c(~input_layer[1065]),
      .d(input_layer[1918]),
      .e(~input_layer[593]),
      .f(input_layer[1761]),
      .y(Y[156]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_94 for neuron157_1
  function_94 neuron157_1 (
      .a(~input_layer[456]),
      .b(input_layer[2168]),
      .c(~input_layer[920]),
      .d(~input_layer[1650]),
      .e(~input_layer[1186]),
      .y(Y[157]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron158_1
  function_10 neuron158_1 (
      .a(input_layer[1662]),
      .b(~input_layer[889]),
      .c(input_layer[1041]),
      .d(~input_layer[872]),
      .y(Y[158]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron159_1
  function_95 neuron159_1 (
      .a(~input_layer[1639]),
      .b(input_layer[1877]),
      .c(~input_layer[1996]),
      .d(input_layer[1743]),
      .y(Y[159]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[160] = 1'b1;

  // instantiate function_26 for neuron161_1
  function_26 neuron161_1 (
      .a(~input_layer[1918]),
      .b(~input_layer[1150]),
      .y(Y[161]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron162_1
  function_24 neuron162_1 (
      .a(~input_layer[832]),
      .y(Y[162]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_96 for neuron163_1
  function_96 neuron163_1 (
      .a(~input_layer[1114]),
      .b(input_layer[1813]),
      .c(input_layer[270]),
      .d(~input_layer[2169]),
      .e(~input_layer[327]),
      .f(~input_layer[2193]),
      .y(Y[163]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron164_1
  function_18 neuron164_1 (
      .a(~input_layer[1277]),
      .b(~input_layer[1191]),
      .c(~input_layer[598]),
      .d(~input_layer[1012]),
      .e(~input_layer[2318]),
      .y(Y[164]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron165_1
  function_54 neuron165_1 (
      .a(input_layer[873]),
      .b(input_layer[1557]),
      .c(input_layer[2066]),
      .d(input_layer[346]),
      .e(input_layer[1869]),
      .f(input_layer[1021]),
      .y(Y[165]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron166_1
  function_18 neuron166_1 (
      .a(~input_layer[1039]),
      .b(~input_layer[1027]),
      .c(~input_layer[2114]),
      .d(~input_layer[1886]),
      .e(~input_layer[2063]),
      .y(Y[166]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron167_1
  function_16 neuron167_1 (
      .a(input_layer[547]),
      .b(input_layer[2237]),
      .c(input_layer[876]),
      .y(Y[167]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron168_1
  function_85 neuron168_1 (
      .a(input_layer[1505]),
      .b(input_layer[776]),
      .c(~input_layer[1203]),
      .d(input_layer[2312]),
      .e(input_layer[1950]),
      .f(~input_layer[1117]),
      .y(Y[168]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron169_1
  function_25 neuron169_1 (
      .a(input_layer[353]),
      .b(input_layer[2151]),
      .c(input_layer[1920]),
      .d(input_layer[1844]),
      .e(input_layer[1061]),
      .y(Y[169]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron170_1
  function_14 neuron170_1 (
      .a(~input_layer[939]),
      .b(~input_layer[2156]),
      .c(~input_layer[1208]),
      .d(input_layer[644]),
      .e(input_layer[637]),
      .y(Y[170]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron171_1
  function_10 neuron171_1 (
      .a(input_layer[1671]),
      .b(input_layer[1622]),
      .c(input_layer[459]),
      .d(~input_layer[1399]),
      .y(Y[171]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron172_1
  function_63 neuron172_1 (
      .a(input_layer[1925]),
      .b(input_layer[1384]),
      .c(input_layer[1828]),
      .d(~input_layer[674]),
      .y(Y[172]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_97 for neuron173_1
  function_97 neuron173_1 (
      .a(input_layer[1070]),
      .b(~input_layer[1671]),
      .c(~input_layer[1991]),
      .d(~input_layer[775]),
      .e(input_layer[151]),
      .f(~input_layer[258]),
      .y(Y[173]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron174_1
  function_0 neuron174_1 (
      .a(~input_layer[1642]),
      .b(input_layer[349]),
      .c(input_layer[2249]),
      .d(input_layer[262]),
      .e(~input_layer[729]),
      .y(Y[174]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_98 for neuron175_1
  function_98 neuron175_1 (
      .a(~input_layer[1612]),
      .b(input_layer[784]),
      .c(input_layer[1276]),
      .d(input_layer[1855]),
      .e(~input_layer[1343]),
      .y(Y[175]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron176_1
  function_54 neuron176_1 (
      .a(input_layer[563]),
      .b(input_layer[1624]),
      .c(input_layer[2312]),
      .d(input_layer[195]),
      .e(input_layer[1721]),
      .f(input_layer[619]),
      .y(Y[176]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron177_1
  function_1 neuron177_1 (
      .a(~input_layer[1421]),
      .b(~input_layer[1253]),
      .c(input_layer[479]),
      .d(~input_layer[1595]),
      .e(~input_layer[2086]),
      .f(~input_layer[2087]),
      .y(Y[177]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron178_1
  function_21 neuron178_1 (
      .a(~input_layer[1382]),
      .b(~input_layer[1828]),
      .c(~input_layer[228]),
      .d(input_layer[1067]),
      .y(Y[178]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron179_1
  function_48 neuron179_1 (
      .a(input_layer[537]),
      .b(input_layer[145]),
      .c(~input_layer[1547]),
      .d(input_layer[2178]),
      .e(~input_layer[148]),
      .y(Y[179]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron180_1
  function_33 neuron180_1 (
      .a(~input_layer[933]),
      .b(~input_layer[1973]),
      .c(~input_layer[1760]),
      .d(input_layer[947]),
      .e(input_layer[949]),
      .y(Y[180]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron181_1
  function_35 neuron181_1 (
      .a(~input_layer[213]),
      .b(input_layer[979]),
      .c(~input_layer[2243]),
      .d(~input_layer[181]),
      .e(input_layer[1022]),
      .y(Y[181]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron182_1
  function_99 neuron182_1 (
      .a(input_layer[1989]),
      .b(input_layer[1811]),
      .c(input_layer[1160]),
      .d(~input_layer[602]),
      .e(input_layer[1561]),
      .f(~input_layer[650]),
      .y(Y[182]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron183_1
  function_67 neuron183_1 (
      .a(input_layer[1333]),
      .b(~input_layer[1665]),
      .c(input_layer[1399]),
      .d(input_layer[2329]),
      .e(~input_layer[556]),
      .y(Y[183]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron184_1
  function_100 neuron184_1 (
      .a(input_layer[1525]),
      .b(~input_layer[1985]),
      .c(input_layer[2301]),
      .y(Y[184]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron185_1
  function_100 neuron185_1 (
      .a(input_layer[1199]),
      .b(~input_layer[1910]),
      .c(~input_layer[934]),
      .y(Y[185]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_101 for neuron186_1
  function_101 neuron186_1 (
      .a(~input_layer[1969]),
      .b(input_layer[1481]),
      .c(~input_layer[1822]),
      .d(input_layer[1486]),
      .e(input_layer[1153]),
      .f(~input_layer[703]),
      .y(Y[186]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron187_1
  function_35 neuron187_1 (
      .a(~input_layer[1971]),
      .b(~input_layer[1356]),
      .c(~input_layer[1991]),
      .d(input_layer[1792]),
      .e(~input_layer[736]),
      .y(Y[187]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_102 for neuron188_1
  function_102 neuron188_1 (
      .a(~input_layer[1479]),
      .b(input_layer[1721]),
      .c(~input_layer[1854]),
      .d(~input_layer[2197]),
      .e(~input_layer[1693]),
      .f(input_layer[2176]),
      .y(Y[188]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_29 for neuron189_1
  function_29 neuron189_1 (
      .a(input_layer[1523]),
      .b(input_layer[225]),
      .c(~input_layer[730]),
      .d(~input_layer[482]),
      .e(~input_layer[699]),
      .f(input_layer[2198]),
      .y(Y[189]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron190_1
  function_35 neuron190_1 (
      .a(~input_layer[1987]),
      .b(~input_layer[1840]),
      .c(~input_layer[755]),
      .d(input_layer[2202]),
      .e(~input_layer[1817]),
      .y(Y[190]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron191_1
  function_10 neuron191_1 (
      .a(~input_layer[1211]),
      .b(input_layer[266]),
      .c(input_layer[1984]),
      .d(input_layer[1511]),
      .y(Y[191]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron192_1
  function_26 neuron192_1 (
      .a(~input_layer[2243]),
      .b(input_layer[1304]),
      .y(Y[192]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron193_1
  function_76 neuron193_1 (
      .a(~input_layer[1469]),
      .b(~input_layer[2244]),
      .c(~input_layer[1113]),
      .d(~input_layer[129]),
      .e(~input_layer[2125]),
      .f(input_layer[1732]),
      .y(Y[193]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_103 for neuron194_1
  function_103 neuron194_1 (
      .a(input_layer[701]),
      .b(input_layer[1449]),
      .c(~input_layer[2152]),
      .d(input_layer[1923]),
      .e(~input_layer[1120]),
      .f(input_layer[2112]),
      .y(Y[194]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron195_1
  function_3 neuron195_1 (
      .a(input_layer[1498]),
      .b(input_layer[669]),
      .c(input_layer[187]),
      .d(input_layer[628]),
      .e(~input_layer[719]),
      .y(Y[195]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron196_1
  function_104 neuron196_1 (
      .a(~input_layer[1896]),
      .b(input_layer[2081]),
      .c(input_layer[195]),
      .y(Y[196]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_105 for neuron197_1
  function_105 neuron197_1 (
      .a(input_layer[992]),
      .b(input_layer[1558]),
      .c(~input_layer[1896]),
      .d(~input_layer[1971]),
      .e(~input_layer[778]),
      .f(input_layer[2054]),
      .y(Y[197]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron198_1
  function_37 neuron198_1 (
      .a(input_layer[765]),
      .b(input_layer[558]),
      .c(~input_layer[1147]),
      .d(input_layer[1987]),
      .e(input_layer[778]),
      .y(Y[198]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_106 for neuron199_1
  function_106 neuron199_1 (
      .a(input_layer[2139]),
      .b(~input_layer[1118]),
      .c(input_layer[1864]),
      .d(~input_layer[2081]),
      .e(input_layer[1649]),
      .f(input_layer[2089]),
      .y(Y[199]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron200_1
  function_16 neuron200_1 (
      .a(input_layer[576]),
      .b(input_layer[538]),
      .c(input_layer[1613]),
      .y(Y[200]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron201_1
  function_107 neuron201_1 (
      .a(~input_layer[1332]),
      .b(input_layer[913]),
      .c(~input_layer[1374]),
      .d(~input_layer[132]),
      .y(Y[201]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron202_1
  function_11 neuron202_1 (
      .a(input_layer[1402]),
      .b(input_layer[2142]),
      .c(input_layer[2008]),
      .d(input_layer[2330]),
      .y(Y[202]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron203_1
  function_10 neuron203_1 (
      .a(input_layer[1607]),
      .b(input_layer[2160]),
      .c(input_layer[447]),
      .d(~input_layer[1415]),
      .y(Y[203]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[204] = 1'b0;

  // instantiate function_108 for neuron205_1
  function_108 neuron205_1 (
      .a(input_layer[1609]),
      .b(~input_layer[1461]),
      .c(~input_layer[1462]),
      .d(~input_layer[1159]),
      .e(input_layer[1697]),
      .f(input_layer[2300]),
      .y(Y[205]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_109 for neuron206_1
  function_109 neuron206_1 (
      .a(input_layer[1754]),
      .b(~input_layer[305]),
      .c(input_layer[2231]),
      .d(input_layer[952]),
      .e(input_layer[1073]),
      .f(input_layer[1788]),
      .y(Y[206]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron207_1
  function_44 neuron207_1 (
      .a(~input_layer[129]),
      .b(~input_layer[2128]),
      .c(input_layer[1784]),
      .y(Y[207]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron208_1
  function_107 neuron208_1 (
      .a(~input_layer[221]),
      .b(input_layer[1333]),
      .c(~input_layer[2310]),
      .d(~input_layer[1092]),
      .y(Y[208]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron209_1
  function_11 neuron209_1 (
      .a(input_layer[2228]),
      .b(input_layer[1757]),
      .c(input_layer[2169]),
      .d(input_layer[2157]),
      .y(Y[209]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron210_1
  function_52 neuron210_1 (
      .a(~input_layer[2217]),
      .b(input_layer[545]),
      .c(~input_layer[1563]),
      .d(input_layer[1715]),
      .e(~input_layer[2237]),
      .y(Y[210]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron211_1
  function_107 neuron211_1 (
      .a(~input_layer[2317]),
      .b(input_layer[2152]),
      .c(~input_layer[300]),
      .d(input_layer[2207]),
      .y(Y[211]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_110 for neuron212_1
  function_110 neuron212_1 (
      .a(~input_layer[434]),
      .b(input_layer[480]),
      .c(input_layer[281]),
      .d(~input_layer[1335]),
      .e(~input_layer[2024]),
      .f(~input_layer[587]),
      .y(Y[212]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron213_1
  function_100 neuron213_1 (
      .a(input_layer[299]),
      .b(~input_layer[1447]),
      .c(input_layer[895]),
      .y(Y[213]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron214_1
  function_67 neuron214_1 (
      .a(input_layer[1991]),
      .b(~input_layer[807]),
      .c(input_layer[1158]),
      .d(input_layer[1151]),
      .e(~input_layer[1957]),
      .y(Y[214]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron215_1
  function_0 neuron215_1 (
      .a(input_layer[1830]),
      .b(input_layer[314]),
      .c(input_layer[1379]),
      .d(input_layer[119]),
      .e(~input_layer[1331]),
      .y(Y[215]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron216_1
  function_0 neuron216_1 (
      .a(input_layer[902]),
      .b(input_layer[1202]),
      .c(input_layer[1278]),
      .d(input_layer[998]),
      .e(input_layer[471]),
      .y(Y[216]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_111 for neuron217_1
  function_111 neuron217_1 (
      .a(input_layer[964]),
      .b(input_layer[1249]),
      .c(input_layer[1074]),
      .d(~input_layer[1216]),
      .e(~input_layer[1353]),
      .f(~input_layer[1488]),
      .y(Y[217]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron218_1
  function_90 neuron218_1 (
      .a(input_layer[1220]),
      .b(~input_layer[276]),
      .c(~input_layer[1641]),
      .d(~input_layer[193]),
      .e(~input_layer[49]),
      .y(Y[218]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron219_1
  function_112 neuron219_1 (
      .a(~input_layer[1189]),
      .b(~input_layer[2027]),
      .c(~input_layer[2042]),
      .d(~input_layer[2224]),
      .e(input_layer[867]),
      .f(~input_layer[1489]),
      .y(Y[219]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron220_1
  function_11 neuron220_1 (
      .a(input_layer[894]),
      .b(input_layer[2160]),
      .c(input_layer[1388]),
      .d(~input_layer[1738]),
      .y(Y[220]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron221_1
  function_113 neuron221_1 (
      .a(input_layer[451]),
      .b(input_layer[1001]),
      .c(~input_layer[553]),
      .d(input_layer[1179]),
      .e(~input_layer[1368]),
      .f(input_layer[1034]),
      .y(Y[221]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron222_1
  function_44 neuron222_1 (
      .a(~input_layer[1784]),
      .b(~input_layer[2216]),
      .c(~input_layer[1941]),
      .y(Y[222]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_114 for neuron223_1
  function_114 neuron223_1 (
      .a(~input_layer[963]),
      .b(~input_layer[1028]),
      .c(input_layer[470]),
      .d(input_layer[1312]),
      .e(~input_layer[1082]),
      .f(input_layer[1893]),
      .y(Y[223]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron224_1
  function_100 neuron224_1 (
      .a(~input_layer[979]),
      .b(~input_layer[1954]),
      .c(input_layer[240]),
      .y(Y[224]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron225_1
  function_42 neuron225_1 (
      .a(input_layer[370]),
      .b(~input_layer[2227]),
      .c(~input_layer[1616]),
      .d(input_layer[1825]),
      .e(input_layer[1184]),
      .y(Y[225]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron226_1
  function_115 neuron226_1 (
      .a(input_layer[1493]),
      .b(~input_layer[372]),
      .c(~input_layer[2005]),
      .d(input_layer[1532]),
      .e(input_layer[365]),
      .y(Y[226]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_114 for neuron227_1
  function_114 neuron227_1 (
      .a(~input_layer[456]),
      .b(input_layer[815]),
      .c(~input_layer[1245]),
      .d(~input_layer[135]),
      .e(input_layer[525]),
      .f(~input_layer[310]),
      .y(Y[227]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron228_1
  function_99 neuron228_1 (
      .a(input_layer[1490]),
      .b(input_layer[1996]),
      .c(input_layer[203]),
      .d(~input_layer[1323]),
      .e(input_layer[1385]),
      .f(~input_layer[651]),
      .y(Y[228]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron229_1
  function_116 neuron229_1 (
      .a(input_layer[1775]),
      .b(~input_layer[1075]),
      .c(~input_layer[1806]),
      .d(input_layer[1679]),
      .y(Y[229]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_81 for neuron230_1
  function_81 neuron230_1 (
      .a(~input_layer[1704]),
      .b(input_layer[1268]),
      .c(~input_layer[2095]),
      .d(input_layer[976]),
      .e(~input_layer[770]),
      .f(~input_layer[1575]),
      .y(Y[230]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron231_1
  function_11 neuron231_1 (
      .a(input_layer[2234]),
      .b(input_layer[774]),
      .c(input_layer[554]),
      .d(input_layer[1874]),
      .y(Y[231]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron232_1
  function_117 neuron232_1 (
      .a(~input_layer[266]),
      .b(input_layer[1308]),
      .c(input_layer[1224]),
      .d(~input_layer[1769]),
      .e(~input_layer[1477]),
      .f(input_layer[2018]),
      .y(Y[232]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_118 for neuron233_1
  function_118 neuron233_1 (
      .a(~input_layer[1284]),
      .b(input_layer[1953]),
      .c(input_layer[1739]),
      .d(input_layer[1024]),
      .e(~input_layer[399]),
      .y(Y[233]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron234_1
  function_119 neuron234_1 (
      .a(input_layer[1870]),
      .b(input_layer[558]),
      .c(input_layer[1791]),
      .d(input_layer[326]),
      .e(input_layer[1982]),
      .f(input_layer[2159]),
      .y(Y[234]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron235_1
  function_12 neuron235_1 (
      .a(~input_layer[299]),
      .b(~input_layer[583]),
      .c(input_layer[1146]),
      .y(Y[235]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron236_1
  function_16 neuron236_1 (
      .a(input_layer[1110]),
      .b(input_layer[574]),
      .c(input_layer[325]),
      .y(Y[236]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron237_1
  function_12 neuron237_1 (
      .a(~input_layer[270]),
      .b(input_layer[1476]),
      .c(~input_layer[1800]),
      .y(Y[237]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron238_1
  function_21 neuron238_1 (
      .a(~input_layer[1408]),
      .b(~input_layer[637]),
      .c(~input_layer[552]),
      .d(~input_layer[1077]),
      .y(Y[238]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron239_1
  function_60 neuron239_1 (
      .a(input_layer[543]),
      .b(~input_layer[121]),
      .c(~input_layer[802]),
      .d(input_layer[1907]),
      .e(~input_layer[149]),
      .f(~input_layer[260]),
      .y(Y[239]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron240_1
  function_76 neuron240_1 (
      .a(~input_layer[1983]),
      .b(~input_layer[1906]),
      .c(~input_layer[1438]),
      .d(~input_layer[1171]),
      .e(~input_layer[546]),
      .f(~input_layer[2178]),
      .y(Y[240]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron241_1
  function_16 neuron241_1 (
      .a(input_layer[1693]),
      .b(input_layer[1959]),
      .c(input_layer[1950]),
      .y(Y[241]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron242_1
  function_26 neuron242_1 (
      .a(~input_layer[1323]),
      .b(~input_layer[1319]),
      .y(Y[242]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron243_1
  function_5 neuron243_1 (
      .a(input_layer[312]),
      .b(input_layer[1142]),
      .y(Y[243]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron244_1
  function_11 neuron244_1 (
      .a(input_layer[518]),
      .b(input_layer[917]),
      .c(input_layer[1582]),
      .d(input_layer[1799]),
      .y(Y[244]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron245_1
  function_120 neuron245_1 (
      .a(input_layer[1075]),
      .b(~input_layer[1783]),
      .c(input_layer[1548]),
      .d(input_layer[1708]),
      .e(input_layer[2285]),
      .f(input_layer[471]),
      .y(Y[245]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_71 for neuron246_1
  function_71 neuron246_1 (
      .a(input_layer[2233]),
      .b(input_layer[498]),
      .c(input_layer[1720]),
      .d(input_layer[869]),
      .e(input_layer[2073]),
      .f(~input_layer[1935]),
      .y(Y[246]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron247_1
  function_121 neuron247_1 (
      .a(~input_layer[1237]),
      .b(input_layer[2329]),
      .c(input_layer[2127]),
      .d(input_layer[187]),
      .e(~input_layer[554]),
      .f(input_layer[1179]),
      .y(Y[247]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron248_1
  function_1 neuron248_1 (
      .a(~input_layer[1577]),
      .b(~input_layer[305]),
      .c(~input_layer[2001]),
      .d(~input_layer[1963]),
      .e(input_layer[974]),
      .f(input_layer[1632]),
      .y(Y[248]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_122 for neuron249_1
  function_122 neuron249_1 (
      .a(input_layer[1167]),
      .b(~input_layer[663]),
      .c(~input_layer[564]),
      .d(~input_layer[566]),
      .e(input_layer[344]),
      .f(input_layer[260]),
      .y(Y[249]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron250_1
  function_35 neuron250_1 (
      .a(~input_layer[2075]),
      .b(~input_layer[826]),
      .c(input_layer[1830]),
      .d(~input_layer[104]),
      .e(~input_layer[396]),
      .y(Y[250]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron251_1
  function_31 neuron251_1 (
      .a(input_layer[1569]),
      .b(input_layer[2130]),
      .c(input_layer[1116]),
      .d(input_layer[1646]),
      .e(input_layer[603]),
      .f(input_layer[1520]),
      .y(Y[251]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron252_1
  function_21 neuron252_1 (
      .a(~input_layer[795]),
      .b(input_layer[373]),
      .c(~input_layer[581]),
      .d(~input_layer[403]),
      .y(Y[252]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron253_1
  function_123 neuron253_1 (
      .a(~input_layer[1502]),
      .b(~input_layer[450]),
      .c(~input_layer[1041]),
      .d(~input_layer[2334]),
      .e(input_layer[843]),
      .f(input_layer[398]),
      .y(Y[253]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron254_1
  function_10 neuron254_1 (
      .a(input_layer[404]),
      .b(input_layer[203]),
      .c(~input_layer[1411]),
      .d(~input_layer[1878]),
      .y(Y[254]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_124 for neuron255_1
  function_124 neuron255_1 (
      .a(~input_layer[956]),
      .b(~input_layer[1124]),
      .c(input_layer[1570]),
      .d(~input_layer[605]),
      .e(~input_layer[1333]),
      .f(~input_layer[146]),
      .y(Y[255]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron256_1
  function_125 neuron256_1 (
      .a(~input_layer[1051]),
      .b(~input_layer[2245]),
      .c(~input_layer[1880]),
      .d(~input_layer[2243]),
      .e(input_layer[1685]),
      .y(Y[256]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron257_1
  function_126 neuron257_1 (
      .a(input_layer[525]),
      .b(input_layer[908]),
      .c(~input_layer[218]),
      .d(~input_layer[954]),
      .e(input_layer[1117]),
      .y(Y[257]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron258_1
  function_25 neuron258_1 (
      .a(input_layer[1492]),
      .b(input_layer[1825]),
      .c(input_layer[1777]),
      .d(input_layer[1674]),
      .e(input_layer[1702]),
      .y(Y[258]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_127 for neuron259_1
  function_127 neuron259_1 (
      .a(input_layer[1986]),
      .b(~input_layer[1735]),
      .c(~input_layer[275]),
      .d(~input_layer[1530]),
      .e(input_layer[674]),
      .f(~input_layer[472]),
      .y(Y[259]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron260_1
  function_128 neuron260_1 (
      .a(input_layer[1133]),
      .b(~input_layer[111]),
      .c(~input_layer[375]),
      .d(~input_layer[1337]),
      .y(Y[260]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron261_1
  function_14 neuron261_1 (
      .a(~input_layer[1418]),
      .b(input_layer[825]),
      .c(~input_layer[1606]),
      .d(~input_layer[2285]),
      .e(~input_layer[1803]),
      .y(Y[261]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron262_1
  function_116 neuron262_1 (
      .a(input_layer[1556]),
      .b(input_layer[1026]),
      .c(~input_layer[434]),
      .d(input_layer[477]),
      .y(Y[262]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_129 for neuron263_1
  function_129 neuron263_1 (
      .a(~input_layer[2230]),
      .b(input_layer[187]),
      .c(input_layer[406]),
      .d(~input_layer[2319]),
      .e(input_layer[866]),
      .f(input_layer[1279]),
      .y(Y[263]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron264_1
  function_18 neuron264_1 (
      .a(~input_layer[1549]),
      .b(~input_layer[744]),
      .c(~input_layer[483]),
      .d(~input_layer[226]),
      .e(~input_layer[318]),
      .y(Y[264]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron265_1
  function_39 neuron265_1 (
      .a(~input_layer[997]),
      .b(~input_layer[1501]),
      .c(input_layer[235]),
      .d(input_layer[1604]),
      .y(Y[265]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron266_1
  function_3 neuron266_1 (
      .a(input_layer[437]),
      .b(input_layer[1438]),
      .c(~input_layer[1466]),
      .d(input_layer[1254]),
      .e(input_layer[1256]),
      .y(Y[266]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron267_1
  function_3 neuron267_1 (
      .a(input_layer[1550]),
      .b(input_layer[2296]),
      .c(~input_layer[1222]),
      .d(input_layer[696]),
      .e(input_layer[2284]),
      .y(Y[267]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron268_1
  function_130 neuron268_1 (
      .a(input_layer[325]),
      .b(~input_layer[1536]),
      .c(input_layer[516]),
      .d(~input_layer[2322]),
      .e(~input_layer[78]),
      .f(input_layer[167]),
      .y(Y[268]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron269_1
  function_131 neuron269_1 (
      .a(input_layer[682]),
      .b(~input_layer[640]),
      .c(~input_layer[1330]),
      .d(~input_layer[2006]),
      .e(input_layer[2336]),
      .f(input_layer[58]),
      .y(Y[269]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron270_1
  function_48 neuron270_1 (
      .a(input_layer[349]),
      .b(~input_layer[549]),
      .c(input_layer[488]),
      .d(input_layer[345]),
      .e(input_layer[919]),
      .y(Y[270]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron271_1
  function_61 neuron271_1 (
      .a(~input_layer[735]),
      .b(~input_layer[2042]),
      .c(input_layer[585]),
      .d(~input_layer[1883]),
      .e(~input_layer[1441]),
      .y(Y[271]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron272_1
  function_131 neuron272_1 (
      .a(~input_layer[1750]),
      .b(~input_layer[1908]),
      .c(input_layer[144]),
      .d(~input_layer[517]),
      .e(~input_layer[1316]),
      .f(~input_layer[331]),
      .y(Y[272]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron273_1
  function_16 neuron273_1 (
      .a(input_layer[641]),
      .b(input_layer[1816]),
      .c(~input_layer[953]),
      .y(Y[273]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron274_1
  function_132 neuron274_1 (
      .a(~input_layer[1727]),
      .b(input_layer[1440]),
      .c(~input_layer[198]),
      .d(~input_layer[1076]),
      .e(input_layer[844]),
      .y(Y[274]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron275_1
  function_24 neuron275_1 (
      .a(~input_layer[1795]),
      .y(Y[275]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron276_1
  function_44 neuron276_1 (
      .a(~input_layer[949]),
      .b(~input_layer[1647]),
      .c(~input_layer[2295]),
      .y(Y[276]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron277_1
  function_63 neuron277_1 (
      .a(input_layer[2034]),
      .b(~input_layer[1232]),
      .c(input_layer[1472]),
      .d(~input_layer[976]),
      .y(Y[277]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron278_1
  function_35 neuron278_1 (
      .a(~input_layer[1367]),
      .b(~input_layer[2143]),
      .c(~input_layer[727]),
      .d(~input_layer[812]),
      .e(input_layer[1783]),
      .y(Y[278]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron279_1
  function_133 neuron279_1 (
      .a(~input_layer[2155]),
      .b(input_layer[1587]),
      .c(input_layer[612]),
      .d(input_layer[828]),
      .e(input_layer[1320]),
      .y(Y[279]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_134 for neuron280_1
  function_134 neuron280_1 (
      .a(input_layer[1410]),
      .b(~input_layer[789]),
      .c(~input_layer[342]),
      .d(input_layer[1093]),
      .e(~input_layer[2137]),
      .f(~input_layer[2072]),
      .y(Y[280]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron281_1
  function_135 neuron281_1 (
      .a(~input_layer[1215]),
      .b(input_layer[2324]),
      .c(input_layer[2311]),
      .d(~input_layer[1382]),
      .e(input_layer[1675]),
      .y(Y[281]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_136 for neuron282_1
  function_136 neuron282_1 (
      .a(~input_layer[1049]),
      .b(~input_layer[2238]),
      .c(input_layer[311]),
      .d(input_layer[1113]),
      .e(~input_layer[853]),
      .f(input_layer[584]),
      .y(Y[282]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron283_1
  function_5 neuron283_1 (
      .a(input_layer[729]),
      .b(input_layer[972]),
      .y(Y[283]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron284_1
  function_113 neuron284_1 (
      .a(input_layer[218]),
      .b(~input_layer[1125]),
      .c(input_layer[112]),
      .d(input_layer[2288]),
      .e(input_layer[694]),
      .f(~input_layer[1263]),
      .y(Y[284]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[285] = 1'b1;

  // instantiate function_137 for neuron286_1
  function_137 neuron286_1 (
      .a(input_layer[1856]),
      .b(input_layer[125]),
      .c(input_layer[887]),
      .d(~input_layer[1205]),
      .e(~input_layer[330]),
      .f(~input_layer[835]),
      .y(Y[286]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_138 for neuron287_1
  function_138 neuron287_1 (
      .a(~input_layer[1030]),
      .b(~input_layer[1124]),
      .c(input_layer[2156]),
      .d(~input_layer[131]),
      .e(input_layer[945]),
      .f(~input_layer[1887]),
      .y(Y[287]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron288_1
  function_107 neuron288_1 (
      .a(~input_layer[1673]),
      .b(~input_layer[233]),
      .c(~input_layer[1501]),
      .d(input_layer[581]),
      .y(Y[288]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron289_1
  function_21 neuron289_1 (
      .a(~input_layer[1569]),
      .b(~input_layer[318]),
      .c(~input_layer[438]),
      .d(~input_layer[2318]),
      .y(Y[289]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron290_1
  function_139 neuron290_1 (
      .a(input_layer[2154]),
      .b(~input_layer[1552]),
      .c(~input_layer[2095]),
      .d(~input_layer[395]),
      .e(~input_layer[319]),
      .y(Y[290]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_140 for neuron291_1
  function_140 neuron291_1 (
      .a(~input_layer[2063]),
      .b(input_layer[858]),
      .c(input_layer[1256]),
      .d(input_layer[1537]),
      .e(~input_layer[1354]),
      .f(~input_layer[1565]),
      .y(Y[291]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_141 for neuron292_1
  function_141 neuron292_1 (
      .a(input_layer[1077]),
      .b(~input_layer[1333]),
      .c(input_layer[2172]),
      .d(input_layer[427]),
      .e(~input_layer[1876]),
      .f(input_layer[2110]),
      .y(Y[292]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_142 for neuron293_1
  function_142 neuron293_1 (
      .a(~input_layer[494]),
      .b(input_layer[1560]),
      .c(~input_layer[1828]),
      .d(input_layer[1025]),
      .e(input_layer[1331]),
      .y(Y[293]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron294_1
  function_21 neuron294_1 (
      .a(~input_layer[711]),
      .b(~input_layer[1632]),
      .c(~input_layer[2213]),
      .d(~input_layer[1951]),
      .y(Y[294]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron295_1
  function_21 neuron295_1 (
      .a(~input_layer[1871]),
      .b(~input_layer[833]),
      .c(input_layer[873]),
      .d(input_layer[780]),
      .y(Y[295]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_121 for neuron296_1
  function_121 neuron296_1 (
      .a(input_layer[958]),
      .b(input_layer[2246]),
      .c(~input_layer[1717]),
      .d(input_layer[1460]),
      .e(input_layer[405]),
      .f(~input_layer[1837]),
      .y(Y[296]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron297_1
  function_14 neuron297_1 (
      .a(~input_layer[908]),
      .b(~input_layer[894]),
      .c(~input_layer[1511]),
      .d(~input_layer[1196]),
      .e(input_layer[786]),
      .y(Y[297]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron298_1
  function_25 neuron298_1 (
      .a(input_layer[850]),
      .b(input_layer[2147]),
      .c(input_layer[1435]),
      .d(input_layer[317]),
      .e(input_layer[2236]),
      .y(Y[298]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_143 for neuron299_1
  function_143 neuron299_1 (
      .a(input_layer[974]),
      .b(input_layer[1423]),
      .c(input_layer[221]),
      .d(~input_layer[625]),
      .e(input_layer[1734]),
      .f(input_layer[629]),
      .y(Y[299]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_144 for neuron300_1
  function_144 neuron300_1 (
      .a(~input_layer[1705]),
      .b(~input_layer[2304]),
      .c(~input_layer[229]),
      .d(input_layer[1526]),
      .e(input_layer[989]),
      .f(~input_layer[783]),
      .y(Y[300]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron301_1
  function_145 neuron301_1 (
      .a(input_layer[765]),
      .b(input_layer[1172]),
      .c(~input_layer[1076]),
      .d(input_layer[1879]),
      .e(input_layer[2050]),
      .f(~input_layer[1035]),
      .y(Y[301]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron302_1
  function_14 neuron302_1 (
      .a(~input_layer[433]),
      .b(~input_layer[1368]),
      .c(~input_layer[2007]),
      .d(~input_layer[1724]),
      .e(~input_layer[943]),
      .y(Y[302]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron303_1
  function_72 neuron303_1 (
      .a(~input_layer[1247]),
      .b(~input_layer[889]),
      .c(~input_layer[453]),
      .d(~input_layer[1432]),
      .e(~input_layer[1747]),
      .y(Y[303]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron304_1
  function_11 neuron304_1 (
      .a(input_layer[816]),
      .b(input_layer[651]),
      .c(input_layer[405]),
      .d(input_layer[2331]),
      .y(Y[304]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron305_1
  function_16 neuron305_1 (
      .a(~input_layer[1041]),
      .b(~input_layer[1389]),
      .c(input_layer[442]),
      .y(Y[305]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron306_1
  function_21 neuron306_1 (
      .a(~input_layer[872]),
      .b(~input_layer[1084]),
      .c(input_layer[1221]),
      .d(input_layer[1609]),
      .y(Y[306]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron307_1
  function_146 neuron307_1 (
      .a(input_layer[1335]),
      .b(input_layer[309]),
      .c(input_layer[657]),
      .d(input_layer[582]),
      .e(~input_layer[563]),
      .y(Y[307]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_147 for neuron308_1
  function_147 neuron308_1 (
      .a(~input_layer[499]),
      .b(input_layer[212]),
      .c(input_layer[210]),
      .d(~input_layer[1614]),
      .e(input_layer[636]),
      .f(~input_layer[1799]),
      .y(Y[308]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron309_1
  function_20 neuron309_1 (
      .a(input_layer[201]),
      .b(~input_layer[1216]),
      .c(input_layer[510]),
      .d(input_layer[2195]),
      .e(input_layer[1937]),
      .f(input_layer[96]),
      .y(Y[309]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron310_1
  function_107 neuron310_1 (
      .a(~input_layer[608]),
      .b(~input_layer[481]),
      .c(input_layer[1136]),
      .d(input_layer[2194]),
      .y(Y[310]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron311_1
  function_11 neuron311_1 (
      .a(input_layer[282]),
      .b(input_layer[441]),
      .c(input_layer[1279]),
      .d(~input_layer[709]),
      .y(Y[311]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron312_1
  function_25 neuron312_1 (
      .a(input_layer[1334]),
      .b(input_layer[681]),
      .c(input_layer[985]),
      .d(input_layer[2245]),
      .e(input_layer[190]),
      .y(Y[312]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[313] = 1'b1;

  // instantiate function_30 for neuron314_1
  function_30 neuron314_1 (
      .a(~input_layer[441]),
      .b(input_layer[148]),
      .c(input_layer[726]),
      .d(input_layer[1920]),
      .y(Y[314]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron315_1
  function_148 neuron315_1 (
      .a(~input_layer[1742]),
      .b(input_layer[775]),
      .c(~input_layer[1732]),
      .d(input_layer[694]),
      .y(Y[315]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron316_1
  function_149 neuron316_1 (
      .a(~input_layer[1246]),
      .b(input_layer[745]),
      .c(~input_layer[1140]),
      .d(input_layer[816]),
      .y(Y[316]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron317_1
  function_107 neuron317_1 (
      .a(~input_layer[2003]),
      .b(~input_layer[284]),
      .c(input_layer[820]),
      .d(input_layer[146]),
      .y(Y[317]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron318_1
  function_3 neuron318_1 (
      .a(input_layer[2215]),
      .b(input_layer[409]),
      .c(input_layer[2292]),
      .d(~input_layer[539]),
      .e(input_layer[1398]),
      .y(Y[318]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron319_1
  function_11 neuron319_1 (
      .a(input_layer[348]),
      .b(input_layer[219]),
      .c(input_layer[274]),
      .d(input_layer[994]),
      .y(Y[319]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron320_1
  function_11 neuron320_1 (
      .a(input_layer[1704]),
      .b(~input_layer[1471]),
      .c(input_layer[2288]),
      .d(input_layer[643]),
      .y(Y[320]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_150 for neuron321_1
  function_150 neuron321_1 (
      .a(input_layer[1627]),
      .b(~input_layer[2146]),
      .c(input_layer[1535]),
      .d(input_layer[187]),
      .e(input_layer[288]),
      .f(input_layer[283]),
      .y(Y[321]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron322_1
  function_67 neuron322_1 (
      .a(input_layer[2230]),
      .b(input_layer[1663]),
      .c(input_layer[2109]),
      .d(input_layer[612]),
      .e(~input_layer[812]),
      .y(Y[322]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron323_1
  function_49 neuron323_1 (
      .a(input_layer[1966]),
      .b(input_layer[139]),
      .c(input_layer[575]),
      .d(input_layer[831]),
      .e(input_layer[1694]),
      .f(input_layer[1351]),
      .y(Y[323]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_151 for neuron324_1
  function_151 neuron324_1 (
      .a(~input_layer[471]),
      .b(input_layer[2064]),
      .c(input_layer[2004]),
      .d(~input_layer[1443]),
      .e(~input_layer[331]),
      .y(Y[324]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron325_1
  function_12 neuron325_1 (
      .a(~input_layer[1899]),
      .b(~input_layer[2203]),
      .c(~input_layer[1874]),
      .y(Y[325]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron326_1
  function_67 neuron326_1 (
      .a(input_layer[1217]),
      .b(input_layer[1833]),
      .c(input_layer[910]),
      .d(input_layer[922]),
      .e(input_layer[1263]),
      .y(Y[326]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron327_1
  function_152 neuron327_1 (
      .a(~input_layer[1170]),
      .b(~input_layer[1729]),
      .c(input_layer[798]),
      .d(~input_layer[1515]),
      .e(input_layer[2227]),
      .f(~input_layer[53]),
      .y(Y[327]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron328_1
  function_26 neuron328_1 (
      .a(input_layer[1124]),
      .b(~input_layer[1422]),
      .y(Y[328]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron329_1
  function_72 neuron329_1 (
      .a(~input_layer[361]),
      .b(~input_layer[1394]),
      .c(input_layer[1809]),
      .d(input_layer[1211]),
      .e(~input_layer[1315]),
      .y(Y[329]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron330_1
  function_25 neuron330_1 (
      .a(input_layer[528]),
      .b(input_layer[2035]),
      .c(input_layer[2318]),
      .d(input_layer[864]),
      .e(input_layer[1427]),
      .y(Y[330]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron331_1
  function_26 neuron331_1 (
      .a(~input_layer[1985]),
      .b(~input_layer[1928]),
      .y(Y[331]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron332_1
  function_24 neuron332_1 (
      .a(~input_layer[1143]),
      .y(Y[332]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron333_1
  function_21 neuron333_1 (
      .a(~input_layer[200]),
      .b(~input_layer[2313]),
      .c(~input_layer[751]),
      .d(~input_layer[1743]),
      .y(Y[333]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron334_1
  function_100 neuron334_1 (
      .a(input_layer[1165]),
      .b(~input_layer[2053]),
      .c(~input_layer[585]),
      .y(Y[334]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_153 for neuron335_1
  function_153 neuron335_1 (
      .a(~input_layer[1301]),
      .b(input_layer[2222]),
      .c(~input_layer[102]),
      .d(~input_layer[2106]),
      .e(~input_layer[1286]),
      .f(~input_layer[80]),
      .y(Y[335]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron336_1
  function_154 neuron336_1 (
      .a(~input_layer[1287]),
      .b(input_layer[1466]),
      .c(input_layer[1900]),
      .d(~input_layer[1489]),
      .e(input_layer[1209]),
      .y(Y[336]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron337_1
  function_155 neuron337_1 (
      .a(input_layer[1052]),
      .b(~input_layer[651]),
      .c(input_layer[130]),
      .d(input_layer[1913]),
      .e(input_layer[756]),
      .y(Y[337]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron338_1
  function_12 neuron338_1 (
      .a(~input_layer[474]),
      .b(~input_layer[765]),
      .c(~input_layer[319]),
      .y(Y[338]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron339_1
  function_21 neuron339_1 (
      .a(~input_layer[971]),
      .b(~input_layer[1713]),
      .c(~input_layer[216]),
      .d(~input_layer[679]),
      .y(Y[339]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron340_1
  function_21 neuron340_1 (
      .a(~input_layer[1625]),
      .b(~input_layer[601]),
      .c(~input_layer[485]),
      .d(~input_layer[452]),
      .y(Y[340]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron341_1
  function_16 neuron341_1 (
      .a(input_layer[1946]),
      .b(input_layer[1924]),
      .c(~input_layer[813]),
      .y(Y[341]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron342_1
  function_125 neuron342_1 (
      .a(~input_layer[534]),
      .b(~input_layer[1813]),
      .c(input_layer[2118]),
      .d(~input_layer[1049]),
      .e(~input_layer[1019]),
      .y(Y[342]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron343_1
  function_40 neuron343_1 (
      .a(~input_layer[1449]),
      .b(~input_layer[653]),
      .c(~input_layer[2240]),
      .d(~input_layer[2214]),
      .e(~input_layer[1272]),
      .f(~input_layer[1671]),
      .y(Y[343]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron344_1
  function_14 neuron344_1 (
      .a(~input_layer[1043]),
      .b(~input_layer[1531]),
      .c(~input_layer[1703]),
      .d(~input_layer[464]),
      .e(input_layer[2330]),
      .y(Y[344]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron345_1
  function_156 neuron345_1 (
      .a(~input_layer[1825]),
      .b(~input_layer[543]),
      .c(input_layer[2198]),
      .d(~input_layer[1961]),
      .e(input_layer[1230]),
      .y(Y[345]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron346_1
  function_21 neuron346_1 (
      .a(~input_layer[448]),
      .b(~input_layer[857]),
      .c(input_layer[1639]),
      .d(~input_layer[951]),
      .y(Y[346]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron347_1
  function_82 neuron347_1 (
      .a(input_layer[190]),
      .b(~input_layer[848]),
      .c(~input_layer[2334]),
      .d(~input_layer[1384]),
      .e(~input_layer[1996]),
      .y(Y[347]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron348_1
  function_3 neuron348_1 (
      .a(input_layer[190]),
      .b(input_layer[2047]),
      .c(~input_layer[1378]),
      .d(~input_layer[440]),
      .e(input_layer[2336]),
      .y(Y[348]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron349_1
  function_67 neuron349_1 (
      .a(input_layer[1606]),
      .b(input_layer[1355]),
      .c(~input_layer[562]),
      .d(input_layer[221]),
      .e(input_layer[566]),
      .y(Y[349]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron350_1
  function_95 neuron350_1 (
      .a(~input_layer[2055]),
      .b(input_layer[132]),
      .c(input_layer[1298]),
      .d(input_layer[634]),
      .y(Y[350]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron351_1
  function_157 neuron351_1 (
      .a(~input_layer[1554]),
      .b(~input_layer[1518]),
      .c(input_layer[543]),
      .d(input_layer[1967]),
      .e(input_layer[1571]),
      .f(input_layer[2255]),
      .y(Y[351]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron352_1
  function_99 neuron352_1 (
      .a(input_layer[933]),
      .b(input_layer[1505]),
      .c(input_layer[613]),
      .d(input_layer[1396]),
      .e(input_layer[411]),
      .f(~input_layer[1569]),
      .y(Y[352]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron353_1
  function_26 neuron353_1 (
      .a(~input_layer[876]),
      .b(~input_layer[1033]),
      .y(Y[353]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron354_1
  function_54 neuron354_1 (
      .a(input_layer[2076]),
      .b(input_layer[1338]),
      .c(~input_layer[1795]),
      .d(input_layer[267]),
      .e(~input_layer[813]),
      .f(~input_layer[1199]),
      .y(Y[354]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_127 for neuron355_1
  function_127 neuron355_1 (
      .a(input_layer[1972]),
      .b(~input_layer[1036]),
      .c(input_layer[1520]),
      .d(input_layer[2070]),
      .e(~input_layer[1571]),
      .f(~input_layer[2181]),
      .y(Y[355]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron356_1
  function_12 neuron356_1 (
      .a(~input_layer[1996]),
      .b(~input_layer[1122]),
      .c(~input_layer[695]),
      .y(Y[356]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron357_1
  function_91 neuron357_1 (
      .a(input_layer[284]),
      .b(input_layer[1255]),
      .c(~input_layer[1134]),
      .d(input_layer[992]),
      .e(~input_layer[1765]),
      .f(~input_layer[1807]),
      .y(Y[357]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_158 for neuron358_1
  function_158 neuron358_1 (
      .a(input_layer[690]),
      .b(input_layer[680]),
      .c(input_layer[2074]),
      .d(~input_layer[228]),
      .e(input_layer[1346]),
      .f(input_layer[106]),
      .y(Y[358]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_159 for neuron359_1
  function_159 neuron359_1 (
      .a(input_layer[953]),
      .b(input_layer[660]),
      .c(input_layer[881]),
      .d(~input_layer[1234]),
      .e(input_layer[1241]),
      .f(input_layer[1589]),
      .y(Y[359]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron360_1
  function_18 neuron360_1 (
      .a(~input_layer[1820]),
      .b(~input_layer[1648]),
      .c(~input_layer[1000]),
      .d(~input_layer[1279]),
      .e(~input_layer[1427]),
      .y(Y[360]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_160 for neuron361_1
  function_160 neuron361_1 (
      .a(input_layer[851]),
      .b(~input_layer[1909]),
      .c(~input_layer[708]),
      .d(input_layer[347]),
      .e(~input_layer[1719]),
      .y(Y[361]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_161 for neuron362_1
  function_161 neuron362_1 (
      .a(~input_layer[315]),
      .b(input_layer[2124]),
      .c(input_layer[2222]),
      .d(~input_layer[305]),
      .e(~input_layer[1656]),
      .f(input_layer[478]),
      .y(Y[362]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron363_1
  function_162 neuron363_1 (
      .a(~input_layer[641]),
      .b(~input_layer[239]),
      .c(~input_layer[861]),
      .d(input_layer[1295]),
      .e(~input_layer[593]),
      .y(Y[363]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron364_1
  function_107 neuron364_1 (
      .a(~input_layer[1239]),
      .b(~input_layer[904]),
      .c(~input_layer[1321]),
      .d(~input_layer[187]),
      .y(Y[364]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron365_1
  function_54 neuron365_1 (
      .a(input_layer[1236]),
      .b(input_layer[2077]),
      .c(input_layer[584]),
      .d(input_layer[1722]),
      .e(input_layer[592]),
      .f(input_layer[1062]),
      .y(Y[365]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_163 for neuron366_1
  function_163 neuron366_1 (
      .a(~input_layer[1227]),
      .b(input_layer[2292]),
      .c(input_layer[1570]),
      .d(~input_layer[443]),
      .e(input_layer[1325]),
      .f(input_layer[44]),
      .y(Y[366]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron367_1
  function_5 neuron367_1 (
      .a(input_layer[1782]),
      .b(~input_layer[1150]),
      .y(Y[367]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron368_1
  function_95 neuron368_1 (
      .a(input_layer[1539]),
      .b(~input_layer[1129]),
      .c(~input_layer[915]),
      .d(input_layer[1053]),
      .y(Y[368]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_164 for neuron369_1
  function_164 neuron369_1 (
      .a(~input_layer[730]),
      .b(input_layer[1468]),
      .c(input_layer[482]),
      .d(~input_layer[2048]),
      .e(~input_layer[2154]),
      .y(Y[369]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron370_1
  function_67 neuron370_1 (
      .a(input_layer[478]),
      .b(input_layer[377]),
      .c(input_layer[1538]),
      .d(~input_layer[609]),
      .e(input_layer[943]),
      .y(Y[370]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron371_1
  function_155 neuron371_1 (
      .a(input_layer[1251]),
      .b(input_layer[1460]),
      .c(input_layer[676]),
      .d(input_layer[1379]),
      .e(~input_layer[1324]),
      .y(Y[371]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron372_1
  function_70 neuron372_1 (
      .a(~input_layer[744]),
      .b(input_layer[1841]),
      .c(~input_layer[1963]),
      .d(~input_layer[672]),
      .e(input_layer[925]),
      .f(input_layer[1559]),
      .y(Y[372]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron373_1
  function_162 neuron373_1 (
      .a(~input_layer[432]),
      .b(input_layer[951]),
      .c(input_layer[293]),
      .d(~input_layer[899]),
      .e(input_layer[1985]),
      .y(Y[373]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron374_1
  function_107 neuron374_1 (
      .a(~input_layer[853]),
      .b(~input_layer[2091]),
      .c(~input_layer[101]),
      .d(~input_layer[1263]),
      .y(Y[374]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron375_1
  function_35 neuron375_1 (
      .a(~input_layer[867]),
      .b(~input_layer[1422]),
      .c(input_layer[1130]),
      .d(~input_layer[1101]),
      .e(~input_layer[438]),
      .y(Y[375]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron376_1
  function_3 neuron376_1 (
      .a(input_layer[2134]),
      .b(input_layer[1676]),
      .c(input_layer[622]),
      .d(input_layer[632]),
      .e(~input_layer[1452]),
      .y(Y[376]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron377_1
  function_26 neuron377_1 (
      .a(~input_layer[1113]),
      .b(~input_layer[2138]),
      .y(Y[377]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron378_1
  function_165 neuron378_1 (
      .a(~input_layer[1451]),
      .b(~input_layer[1842]),
      .c(input_layer[965]),
      .d(input_layer[1967]),
      .e(~input_layer[840]),
      .f(input_layer[2107]),
      .y(Y[378]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron379_1
  function_107 neuron379_1 (
      .a(~input_layer[902]),
      .b(~input_layer[2315]),
      .c(~input_layer[1397]),
      .d(~input_layer[1070]),
      .y(Y[379]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron380_1
  function_3 neuron380_1 (
      .a(input_layer[540]),
      .b(input_layer[947]),
      .c(input_layer[1144]),
      .d(input_layer[544]),
      .e(input_layer[2022]),
      .y(Y[380]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron381_1
  function_104 neuron381_1 (
      .a(input_layer[1841]),
      .b(~input_layer[306]),
      .c(~input_layer[1300]),
      .y(Y[381]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron382_1
  function_3 neuron382_1 (
      .a(input_layer[747]),
      .b(input_layer[116]),
      .c(input_layer[1045]),
      .d(input_layer[566]),
      .e(input_layer[594]),
      .y(Y[382]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron383_1
  function_149 neuron383_1 (
      .a(~input_layer[980]),
      .b(~input_layer[591]),
      .c(~input_layer[126]),
      .d(input_layer[1977]),
      .y(Y[383]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_7 for neuron384_1
  function_7 neuron384_1 (
      .a(input_layer[896]),
      .b(input_layer[676]),
      .c(~input_layer[2240]),
      .d(~input_layer[1677]),
      .e(input_layer[2016]),
      .f(~input_layer[2340]),
      .y(Y[384]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron385_1
  function_24 neuron385_1 (
      .a(~input_layer[886]),
      .y(Y[385]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron386_1
  function_3 neuron386_1 (
      .a(input_layer[1605]),
      .b(input_layer[530]),
      .c(~input_layer[1381]),
      .d(~input_layer[1136]),
      .e(input_layer[775]),
      .y(Y[386]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron387_1
  function_11 neuron387_1 (
      .a(input_layer[1103]),
      .b(input_layer[2057]),
      .c(input_layer[1979]),
      .d(input_layer[1433]),
      .y(Y[387]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron388_1
  function_65 neuron388_1 (
      .a(~input_layer[559]),
      .b(~input_layer[2136]),
      .c(~input_layer[2090]),
      .d(input_layer[985]),
      .e(~input_layer[1676]),
      .f(input_layer[111]),
      .y(Y[388]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_166 for neuron389_1
  function_166 neuron389_1 (
      .a(~input_layer[275]),
      .b(~input_layer[121]),
      .c(input_layer[978]),
      .d(input_layer[671]),
      .e(input_layer[677]),
      .f(~input_layer[552]),
      .y(Y[389]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron390_1
  function_5 neuron390_1 (
      .a(~input_layer[736]),
      .b(input_layer[2242]),
      .y(Y[390]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron391_1
  function_37 neuron391_1 (
      .a(input_layer[1278]),
      .b(~input_layer[1419]),
      .c(~input_layer[1798]),
      .d(input_layer[760]),
      .e(~input_layer[1642]),
      .y(Y[391]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron392_1
  function_167 neuron392_1 (
      .a(~input_layer[2170]),
      .b(~input_layer[1054]),
      .c(input_layer[1548]),
      .d(input_layer[695]),
      .e(input_layer[2287]),
      .y(Y[392]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_168 for neuron393_1
  function_168 neuron393_1 (
      .a(~input_layer[770]),
      .b(input_layer[965]),
      .c(~input_layer[1483]),
      .d(input_layer[940]),
      .e(~input_layer[697]),
      .f(~input_layer[1514]),
      .y(Y[393]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron394_1
  function_67 neuron394_1 (
      .a(input_layer[790]),
      .b(input_layer[2320]),
      .c(~input_layer[1651]),
      .d(input_layer[549]),
      .e(~input_layer[1248]),
      .y(Y[394]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron395_1
  function_169 neuron395_1 (
      .a(input_layer[278]),
      .b(~input_layer[1629]),
      .c(input_layer[386]),
      .d(input_layer[1787]),
      .e(input_layer[2281]),
      .f(input_layer[2068]),
      .y(Y[395]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron396_1
  function_154 neuron396_1 (
      .a(input_layer[583]),
      .b(input_layer[490]),
      .c(~input_layer[2127]),
      .d(~input_layer[2131]),
      .e(input_layer[1458]),
      .y(Y[396]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron397_1
  function_170 neuron397_1 (
      .a(~input_layer[110]),
      .b(~input_layer[118]),
      .c(input_layer[979]),
      .d(~input_layer[1378]),
      .e(~input_layer[179]),
      .y(Y[397]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron398_1
  function_72 neuron398_1 (
      .a(input_layer[570]),
      .b(~input_layer[2218]),
      .c(~input_layer[191]),
      .d(~input_layer[2332]),
      .e(input_layer[1850]),
      .y(Y[398]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_171 for neuron399_1
  function_171 neuron399_1 (
      .a(input_layer[1819]),
      .b(~input_layer[143]),
      .c(~input_layer[344]),
      .d(input_layer[820]),
      .e(~input_layer[358]),
      .f(~input_layer[266]),
      .y(Y[399]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron400_1
  function_148 neuron400_1 (
      .a(~input_layer[1997]),
      .b(input_layer[2112]),
      .c(input_layer[1062]),
      .d(~input_layer[1529]),
      .y(Y[400]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron401_1
  function_16 neuron401_1 (
      .a(~input_layer[1141]),
      .b(input_layer[329]),
      .c(input_layer[96]),
      .y(Y[401]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron402_1
  function_26 neuron402_1 (
      .a(input_layer[902]),
      .b(~input_layer[1352]),
      .y(Y[402]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron403_1
  function_90 neuron403_1 (
      .a(~input_layer[1462]),
      .b(~input_layer[439]),
      .c(input_layer[490]),
      .d(~input_layer[1348]),
      .e(~input_layer[969]),
      .y(Y[403]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron404_1
  function_18 neuron404_1 (
      .a(~input_layer[451]),
      .b(~input_layer[613]),
      .c(input_layer[312]),
      .d(~input_layer[2199]),
      .e(~input_layer[1844]),
      .y(Y[404]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron405_1
  function_14 neuron405_1 (
      .a(~input_layer[1700]),
      .b(~input_layer[304]),
      .c(~input_layer[1630]),
      .d(~input_layer[1436]),
      .e(input_layer[814]),
      .y(Y[405]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron406_1
  function_0 neuron406_1 (
      .a(input_layer[374]),
      .b(~input_layer[550]),
      .c(input_layer[2023]),
      .d(input_layer[1258]),
      .e(input_layer[1061]),
      .y(Y[406]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron407_1
  function_3 neuron407_1 (
      .a(input_layer[1158]),
      .b(input_layer[1586]),
      .c(input_layer[1327]),
      .d(input_layer[209]),
      .e(input_layer[1926]),
      .y(Y[407]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron408_1
  function_3 neuron408_1 (
      .a(input_layer[386]),
      .b(input_layer[396]),
      .c(input_layer[284]),
      .d(input_layer[1219]),
      .e(input_layer[98]),
      .y(Y[408]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron409_1
  function_100 neuron409_1 (
      .a(input_layer[2229]),
      .b(input_layer[928]),
      .c(~input_layer[1687]),
      .y(Y[409]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron410_1
  function_10 neuron410_1 (
      .a(input_layer[1463]),
      .b(input_layer[849]),
      .c(input_layer[1946]),
      .d(~input_layer[1124]),
      .y(Y[410]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron411_1
  function_17 neuron411_1 (
      .a(~input_layer[908]),
      .b(input_layer[1695]),
      .c(~input_layer[1182]),
      .d(~input_layer[2244]),
      .e(~input_layer[1712]),
      .f(input_layer[2007]),
      .y(Y[411]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron412_1
  function_172 neuron412_1 (
      .a(~input_layer[1690]),
      .b(~input_layer[1521]),
      .c(~input_layer[963]),
      .d(input_layer[2165]),
      .e(input_layer[265]),
      .f(~input_layer[443]),
      .y(Y[412]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_173 for neuron413_1
  function_173 neuron413_1 (
      .a(~input_layer[739]),
      .b(input_layer[719]),
      .c(input_layer[1927]),
      .d(~input_layer[787]),
      .e(input_layer[1855]),
      .f(~input_layer[2067]),
      .y(Y[413]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron414_1
  function_3 neuron414_1 (
      .a(input_layer[810]),
      .b(input_layer[2205]),
      .c(input_layer[1925]),
      .d(input_layer[480]),
      .e(~input_layer[1048]),
      .y(Y[414]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron415_1
  function_10 neuron415_1 (
      .a(input_layer[1338]),
      .b(input_layer[1114]),
      .c(~input_layer[368]),
      .d(input_layer[326]),
      .y(Y[415]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron416_1
  function_116 neuron416_1 (
      .a(input_layer[1663]),
      .b(input_layer[1519]),
      .c(~input_layer[676]),
      .d(input_layer[1651]),
      .y(Y[416]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron417_1
  function_42 neuron417_1 (
      .a(input_layer[353]),
      .b(input_layer[891]),
      .c(~input_layer[794]),
      .d(input_layer[1974]),
      .e(input_layer[98]),
      .y(Y[417]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron418_1
  function_93 neuron418_1 (
      .a(~input_layer[1786]),
      .b(~input_layer[195]),
      .c(input_layer[1310]),
      .d(~input_layer[639]),
      .e(input_layer[2067]),
      .f(~input_layer[1345]),
      .y(Y[418]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron419_1
  function_25 neuron419_1 (
      .a(input_layer[1779]),
      .b(input_layer[1052]),
      .c(input_layer[209]),
      .d(input_layer[1437]),
      .e(input_layer[1625]),
      .y(Y[419]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron420_1
  function_5 neuron420_1 (
      .a(~input_layer[1373]),
      .b(input_layer[348]),
      .y(Y[420]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron421_1
  function_12 neuron421_1 (
      .a(~input_layer[2218]),
      .b(input_layer[472]),
      .c(input_layer[1057]),
      .y(Y[421]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron422_1
  function_25 neuron422_1 (
      .a(input_layer[1336]),
      .b(input_layer[298]),
      .c(input_layer[289]),
      .d(~input_layer[576]),
      .e(input_layer[2083]),
      .y(Y[422]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron423_1
  function_21 neuron423_1 (
      .a(~input_layer[2047]),
      .b(~input_layer[2152]),
      .c(input_layer[1725]),
      .d(~input_layer[1020]),
      .y(Y[423]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron424_1
  function_17 neuron424_1 (
      .a(~input_layer[283]),
      .b(input_layer[1056]),
      .c(~input_layer[1633]),
      .d(~input_layer[1299]),
      .e(~input_layer[1178]),
      .f(~input_layer[1]),
      .y(Y[424]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_174 for neuron425_1
  function_174 neuron425_1 (
      .a(~input_layer[224]),
      .b(input_layer[1651]),
      .c(input_layer[1350]),
      .d(input_layer[1714]),
      .e(input_layer[643]),
      .f(~input_layer[2153]),
      .y(Y[425]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron426_1
  function_175 neuron426_1 (
      .a(~input_layer[2211]),
      .b(input_layer[788]),
      .c(~input_layer[829]),
      .d(~input_layer[1974]),
      .e(input_layer[1938]),
      .y(Y[426]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron427_1
  function_18 neuron427_1 (
      .a(~input_layer[1861]),
      .b(~input_layer[1698]),
      .c(~input_layer[1662]),
      .d(~input_layer[1657]),
      .e(~input_layer[300]),
      .y(Y[427]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron428_1
  function_116 neuron428_1 (
      .a(input_layer[2119]),
      .b(input_layer[798]),
      .c(~input_layer[903]),
      .d(input_layer[448]),
      .y(Y[428]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_176 for neuron429_1
  function_176 neuron429_1 (
      .a(input_layer[202]),
      .b(input_layer[1373]),
      .c(input_layer[473]),
      .d(~input_layer[703]),
      .e(~input_layer[2297]),
      .f(~input_layer[711]),
      .y(Y[429]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron430_1
  function_25 neuron430_1 (
      .a(input_layer[1362]),
      .b(~input_layer[1814]),
      .c(input_layer[1162]),
      .d(input_layer[2071]),
      .e(input_layer[2324]),
      .y(Y[430]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron431_1
  function_1 neuron431_1 (
      .a(~input_layer[362]),
      .b(~input_layer[1352]),
      .c(input_layer[982]),
      .d(~input_layer[1803]),
      .e(~input_layer[1280]),
      .f(~input_layer[1548]),
      .y(Y[431]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron432_1
  function_21 neuron432_1 (
      .a(~input_layer[1712]),
      .b(~input_layer[214]),
      .c(~input_layer[553]),
      .d(input_layer[1557]),
      .y(Y[432]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron433_1
  function_67 neuron433_1 (
      .a(input_layer[206]),
      .b(input_layer[1074]),
      .c(input_layer[301]),
      .d(~input_layer[1659]),
      .e(input_layer[1718]),
      .y(Y[433]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_177 for neuron434_1
  function_177 neuron434_1 (
      .a(input_layer[2118]),
      .b(~input_layer[991]),
      .c(~input_layer[105]),
      .d(input_layer[478]),
      .e(~input_layer[838]),
      .f(~input_layer[2142]),
      .y(Y[434]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron435_1
  function_113 neuron435_1 (
      .a(input_layer[631]),
      .b(input_layer[1617]),
      .c(input_layer[965]),
      .d(~input_layer[1313]),
      .e(input_layer[2325]),
      .f(input_layer[672]),
      .y(Y[435]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron436_1
  function_28 neuron436_1 (
      .a(input_layer[808]),
      .b(input_layer[2035]),
      .c(~input_layer[1552]),
      .d(input_layer[700]),
      .e(~input_layer[640]),
      .f(input_layer[1393]),
      .y(Y[436]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron437_1
  function_157 neuron437_1 (
      .a(~input_layer[1653]),
      .b(~input_layer[401]),
      .c(~input_layer[1044]),
      .d(input_layer[1185]),
      .e(input_layer[238]),
      .f(~input_layer[110]),
      .y(Y[437]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_178 for neuron438_1
  function_178 neuron438_1 (
      .a(~input_layer[1017]),
      .b(~input_layer[1087]),
      .c(~input_layer[1055]),
      .d(input_layer[1046]),
      .e(input_layer[300]),
      .f(input_layer[144]),
      .y(Y[438]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron439_1
  function_1 neuron439_1 (
      .a(~input_layer[1714]),
      .b(~input_layer[439]),
      .c(~input_layer[493]),
      .d(~input_layer[1593]),
      .e(input_layer[816]),
      .f(input_layer[1395]),
      .y(Y[439]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron440_1
  function_179 neuron440_1 (
      .a(input_layer[884]),
      .b(input_layer[1605]),
      .c(~input_layer[129]),
      .d(~input_layer[1253]),
      .e(~input_layer[1921]),
      .y(Y[440]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron441_1
  function_139 neuron441_1 (
      .a(input_layer[851]),
      .b(~input_layer[468]),
      .c(~input_layer[1725]),
      .d(~input_layer[1715]),
      .e(input_layer[47]),
      .y(Y[441]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron442_1
  function_67 neuron442_1 (
      .a(input_layer[213]),
      .b(input_layer[1465]),
      .c(~input_layer[1620]),
      .d(~input_layer[1485]),
      .e(input_layer[130]),
      .y(Y[442]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron443_1
  function_11 neuron443_1 (
      .a(input_layer[638]),
      .b(input_layer[1604]),
      .c(input_layer[1943]),
      .d(input_layer[1028]),
      .y(Y[443]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron444_1
  function_92 neuron444_1 (
      .a(~input_layer[305]),
      .b(input_layer[491]),
      .c(input_layer[2304]),
      .d(~input_layer[2044]),
      .y(Y[444]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron445_1
  function_14 neuron445_1 (
      .a(~input_layer[863]),
      .b(~input_layer[2147]),
      .c(~input_layer[2203]),
      .d(~input_layer[1724]),
      .e(input_layer[2091]),
      .y(Y[445]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron446_1
  function_14 neuron446_1 (
      .a(~input_layer[1667]),
      .b(~input_layer[492]),
      .c(~input_layer[1584]),
      .d(input_layer[1868]),
      .e(input_layer[1940]),
      .y(Y[446]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron447_1
  function_8 neuron447_1 (
      .a(~input_layer[319]),
      .b(~input_layer[1172]),
      .c(input_layer[1648]),
      .d(input_layer[996]),
      .e(input_layer[1615]),
      .f(~input_layer[153]),
      .y(Y[447]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_180 for neuron448_1
  function_180 neuron448_1 (
      .a(input_layer[551]),
      .b(~input_layer[952]),
      .c(~input_layer[863]),
      .d(input_layer[890]),
      .e(~input_layer[724]),
      .y(Y[448]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron449_1
  function_116 neuron449_1 (
      .a(input_layer[1667]),
      .b(input_layer[1708]),
      .c(input_layer[470]),
      .d(input_layer[1394]),
      .y(Y[449]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron450_1
  function_63 neuron450_1 (
      .a(input_layer[209]),
      .b(input_layer[1557]),
      .c(~input_layer[935]),
      .d(input_layer[143]),
      .y(Y[450]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron451_1
  function_125 neuron451_1 (
      .a(input_layer[1887]),
      .b(~input_layer[2321]),
      .c(~input_layer[369]),
      .d(input_layer[1055]),
      .e(input_layer[733]),
      .y(Y[451]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron452_1
  function_181 neuron452_1 (
      .a(~input_layer[1839]),
      .b(~input_layer[1373]),
      .c(~input_layer[822]),
      .d(input_layer[1873]),
      .e(~input_layer[925]),
      .f(~input_layer[1281]),
      .y(Y[452]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron453_1
  function_14 neuron453_1 (
      .a(~input_layer[1410]),
      .b(~input_layer[469]),
      .c(~input_layer[1070]),
      .d(input_layer[714]),
      .e(~input_layer[1342]),
      .y(Y[453]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_182 for neuron454_1
  function_182 neuron454_1 (
      .a(input_layer[1201]),
      .b(~input_layer[738]),
      .c(input_layer[331]),
      .d(~input_layer[1076]),
      .e(input_layer[178]),
      .f(input_layer[704]),
      .y(Y[454]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron455_1
  function_183 neuron455_1 (
      .a(input_layer[284]),
      .b(~input_layer[1858]),
      .c(input_layer[709]),
      .d(input_layer[987]),
      .e(~input_layer[1229]),
      .f(~input_layer[445]),
      .y(Y[455]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron456_1
  function_76 neuron456_1 (
      .a(~input_layer[770]),
      .b(~input_layer[2234]),
      .c(~input_layer[2297]),
      .d(input_layer[1386]),
      .e(~input_layer[546]),
      .f(input_layer[282]),
      .y(Y[456]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron457_1
  function_11 neuron457_1 (
      .a(input_layer[1291]),
      .b(input_layer[1586]),
      .c(input_layer[750]),
      .d(input_layer[649]),
      .y(Y[457]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_184 for neuron458_1
  function_184 neuron458_1 (
      .a(~input_layer[299]),
      .b(~input_layer[854]),
      .c(input_layer[1100]),
      .d(input_layer[1273]),
      .e(~input_layer[1568]),
      .y(Y[458]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron459_1
  function_149 neuron459_1 (
      .a(~input_layer[1825]),
      .b(input_layer[1566]),
      .c(~input_layer[1087]),
      .d(input_layer[240]),
      .y(Y[459]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron460_1
  function_21 neuron460_1 (
      .a(~input_layer[1875]),
      .b(~input_layer[2005]),
      .c(~input_layer[2220]),
      .d(input_layer[1547]),
      .y(Y[460]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_185 for neuron461_1
  function_185 neuron461_1 (
      .a(input_layer[412]),
      .b(~input_layer[1872]),
      .c(input_layer[134]),
      .d(input_layer[569]),
      .e(~input_layer[374]),
      .f(input_layer[242]),
      .y(Y[461]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_186 for neuron462_1
  function_186 neuron462_1 (
      .a(~input_layer[1524]),
      .b(input_layer[2200]),
      .c(input_layer[128]),
      .d(input_layer[635]),
      .e(input_layer[835]),
      .f(input_layer[550]),
      .y(Y[462]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron463_1
  function_76 neuron463_1 (
      .a(~input_layer[1584]),
      .b(~input_layer[356]),
      .c(input_layer[1138]),
      .d(~input_layer[234]),
      .e(~input_layer[2027]),
      .f(input_layer[2164]),
      .y(Y[463]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron464_1
  function_18 neuron464_1 (
      .a(~input_layer[1734]),
      .b(~input_layer[1491]),
      .c(~input_layer[1838]),
      .d(~input_layer[1922]),
      .e(~input_layer[685]),
      .y(Y[464]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_187 for neuron465_1
  function_187 neuron465_1 (
      .a(input_layer[1070]),
      .b(input_layer[2213]),
      .c(~input_layer[661]),
      .d(~input_layer[1451]),
      .e(input_layer[1463]),
      .f(input_layer[817]),
      .y(Y[465]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_171 for neuron466_1
  function_171 neuron466_1 (
      .a(~input_layer[1045]),
      .b(input_layer[1061]),
      .c(input_layer[2329]),
      .d(~input_layer[371]),
      .e(input_layer[958]),
      .f(~input_layer[2148]),
      .y(Y[466]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron467_1
  function_188 neuron467_1 (
      .a(input_layer[642]),
      .b(~input_layer[1729]),
      .c(input_layer[675]),
      .d(input_layer[376]),
      .e(input_layer[2342]),
      .f(~input_layer[9]),
      .y(Y[467]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron468_1
  function_16 neuron468_1 (
      .a(input_layer[970]),
      .b(input_layer[282]),
      .c(input_layer[363]),
      .y(Y[468]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron469_1
  function_67 neuron469_1 (
      .a(input_layer[1584]),
      .b(~input_layer[798]),
      .c(input_layer[1452]),
      .d(input_layer[1258]),
      .e(~input_layer[1638]),
      .y(Y[469]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron470_1
  function_5 neuron470_1 (
      .a(input_layer[553]),
      .b(~input_layer[371]),
      .y(Y[470]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_189 for neuron471_1
  function_189 neuron471_1 (
      .a(~input_layer[1791]),
      .b(input_layer[434]),
      .c(~input_layer[150]),
      .d(input_layer[733]),
      .e(input_layer[1929]),
      .y(Y[471]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[472] = 1'b0;

  // instantiate function_48 for neuron473_1
  function_48 neuron473_1 (
      .a(input_layer[887]),
      .b(input_layer[202]),
      .c(~input_layer[1239]),
      .d(input_layer[2066]),
      .e(input_layer[1920]),
      .y(Y[473]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_190 for neuron474_1
  function_190 neuron474_1 (
      .a(~input_layer[961]),
      .b(input_layer[2210]),
      .c(~input_layer[366]),
      .d(input_layer[2286]),
      .e(~input_layer[2046]),
      .f(input_layer[1061]),
      .y(Y[474]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron475_1
  function_18 neuron475_1 (
      .a(~input_layer[1893]),
      .b(~input_layer[2289]),
      .c(~input_layer[2111]),
      .d(~input_layer[245]),
      .e(~input_layer[2079]),
      .y(Y[475]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron476_1
  function_3 neuron476_1 (
      .a(input_layer[1628]),
      .b(input_layer[295]),
      .c(input_layer[496]),
      .d(~input_layer[1155]),
      .e(input_layer[1441]),
      .y(Y[476]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_191 for neuron477_1
  function_191 neuron477_1 (
      .a(input_layer[2036]),
      .b(input_layer[1018]),
      .c(input_layer[500]),
      .d(~input_layer[1253]),
      .e(input_layer[1268]),
      .f(~input_layer[457]),
      .y(Y[477]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron478_1
  function_192 neuron478_1 (
      .a(~input_layer[1782]),
      .b(~input_layer[1945]),
      .c(~input_layer[1778]),
      .d(~input_layer[414]),
      .e(input_layer[2305]),
      .f(input_layer[948]),
      .y(Y[478]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron479_1
  function_5 neuron479_1 (
      .a(input_layer[1281]),
      .b(input_layer[509]),
      .y(Y[479]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron480_1
  function_12 neuron480_1 (
      .a(~input_layer[2062]),
      .b(input_layer[723]),
      .c(~input_layer[2325]),
      .y(Y[480]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron481_1
  function_193 neuron481_1 (
      .a(input_layer[1032]),
      .b(input_layer[752]),
      .c(~input_layer[1438]),
      .d(input_layer[571]),
      .e(~input_layer[1653]),
      .f(input_layer[705]),
      .y(Y[481]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[482] = 1'b1;

  // instantiate function_194 for neuron483_1
  function_194 neuron483_1 (
      .a(input_layer[1791]),
      .b(~input_layer[1377]),
      .c(~input_layer[488]),
      .d(input_layer[229]),
      .e(~input_layer[2167]),
      .f(input_layer[973]),
      .y(Y[483]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron484_1
  function_156 neuron484_1 (
      .a(~input_layer[1132]),
      .b(input_layer[1415]),
      .c(input_layer[1390]),
      .d(~input_layer[1875]),
      .e(input_layer[646]),
      .y(Y[484]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron485_1
  function_11 neuron485_1 (
      .a(input_layer[1066]),
      .b(input_layer[993]),
      .c(input_layer[382]),
      .d(~input_layer[738]),
      .y(Y[485]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron486_1
  function_115 neuron486_1 (
      .a(input_layer[2116]),
      .b(input_layer[483]),
      .c(input_layer[1435]),
      .d(~input_layer[2312]),
      .e(~input_layer[714]),
      .y(Y[486]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron487_1
  function_24 neuron487_1 (
      .a(~input_layer[1611]),
      .y(Y[487]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron488_1
  function_195 neuron488_1 (
      .a(input_layer[743]),
      .b(input_layer[849]),
      .c(~input_layer[1486]),
      .d(~input_layer[2082]),
      .e(input_layer[566]),
      .f(input_layer[1596]),
      .y(Y[488]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron489_1
  function_16 neuron489_1 (
      .a(input_layer[1529]),
      .b(input_layer[1255]),
      .c(~input_layer[1213]),
      .y(Y[489]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron490_1
  function_26 neuron490_1 (
      .a(~input_layer[1907]),
      .b(~input_layer[1256]),
      .y(Y[490]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron491_1
  function_67 neuron491_1 (
      .a(input_layer[1870]),
      .b(input_layer[295]),
      .c(input_layer[2118]),
      .d(input_layer[1167]),
      .e(~input_layer[2072]),
      .y(Y[491]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_196 for neuron492_1
  function_196 neuron492_1 (
      .a(~input_layer[813]),
      .b(input_layer[137]),
      .c(input_layer[497]),
      .d(input_layer[151]),
      .e(input_layer[2093]),
      .f(input_layer[1431]),
      .y(Y[492]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron493_1
  function_107 neuron493_1 (
      .a(~input_layer[1713]),
      .b(~input_layer[2300]),
      .c(input_layer[1560]),
      .d(~input_layer[229]),
      .y(Y[493]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron494_1
  function_25 neuron494_1 (
      .a(input_layer[2312]),
      .b(~input_layer[1107]),
      .c(input_layer[678]),
      .d(input_layer[2288]),
      .e(input_layer[135]),
      .y(Y[494]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_197 for neuron495_1
  function_197 neuron495_1 (
      .a(input_layer[223]),
      .b(~input_layer[2219]),
      .c(~input_layer[1245]),
      .d(input_layer[532]),
      .e(~input_layer[1963]),
      .f(input_layer[1193]),
      .y(Y[495]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron496_1
  function_89 neuron496_1 (
      .a(input_layer[2121]),
      .b(input_layer[2245]),
      .c(~input_layer[684]),
      .d(input_layer[2135]),
      .e(input_layer[1488]),
      .f(input_layer[214]),
      .y(Y[496]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron497_1
  function_21 neuron497_1 (
      .a(~input_layer[1691]),
      .b(~input_layer[2203]),
      .c(~input_layer[1972]),
      .d(input_layer[183]),
      .y(Y[497]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron498_1
  function_48 neuron498_1 (
      .a(input_layer[2075]),
      .b(~input_layer[1734]),
      .c(input_layer[1336]),
      .d(input_layer[1892]),
      .e(~input_layer[396]),
      .y(Y[498]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron499_1
  function_12 neuron499_1 (
      .a(~input_layer[878]),
      .b(input_layer[1402]),
      .c(~input_layer[486]),
      .y(Y[499]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_198 for neuron500_1
  function_198 neuron500_1 (
      .a(input_layer[656]),
      .b(input_layer[1000]),
      .c(~input_layer[2249]),
      .d(~input_layer[1113]),
      .e(input_layer[536]),
      .y(Y[500]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_199 for neuron501_1
  function_199 neuron501_1 (
      .a(~input_layer[608]),
      .b(input_layer[1828]),
      .c(input_layer[487]),
      .d(~input_layer[1946]),
      .e(input_layer[1292]),
      .f(~input_layer[692]),
      .y(Y[501]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron502_1
  function_170 neuron502_1 (
      .a(~input_layer[521]),
      .b(~input_layer[528]),
      .c(input_layer[1072]),
      .d(~input_layer[1363]),
      .e(input_layer[1349]),
      .y(Y[502]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_200 for neuron503_1
  function_200 neuron503_1 (
      .a(input_layer[1629]),
      .b(~input_layer[2028]),
      .c(input_layer[262]),
      .d(input_layer[418]),
      .e(~input_layer[248]),
      .f(input_layer[1]),
      .y(Y[503]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_127 for neuron504_1
  function_127 neuron504_1 (
      .a(input_layer[2087]),
      .b(~input_layer[1443]),
      .c(~input_layer[549]),
      .d(~input_layer[603]),
      .e(input_layer[896]),
      .f(~input_layer[1869]),
      .y(Y[504]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron505_1
  function_95 neuron505_1 (
      .a(~input_layer[401]),
      .b(input_layer[698]),
      .c(input_layer[775]),
      .d(~input_layer[1490]),
      .y(Y[505]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron506_1
  function_21 neuron506_1 (
      .a(~input_layer[368]),
      .b(~input_layer[745]),
      .c(~input_layer[832]),
      .d(~input_layer[1679]),
      .y(Y[506]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron507_1
  function_45 neuron507_1 (
      .a(~input_layer[1402]),
      .b(~input_layer[531]),
      .c(~input_layer[696]),
      .d(~input_layer[441]),
      .e(~input_layer[1097]),
      .f(input_layer[2046]),
      .y(Y[507]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_201 for neuron508_1
  function_201 neuron508_1 (
      .a(input_layer[1049]),
      .b(input_layer[958]),
      .c(~input_layer[1401]),
      .d(~input_layer[2334]),
      .e(~input_layer[22]),
      .y(Y[508]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron509_1
  function_116 neuron509_1 (
      .a(input_layer[1053]),
      .b(~input_layer[1447]),
      .c(input_layer[1675]),
      .d(input_layer[107]),
      .y(Y[509]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron510_1
  function_90 neuron510_1 (
      .a(~input_layer[1578]),
      .b(~input_layer[450]),
      .c(~input_layer[1707]),
      .d(~input_layer[777]),
      .e(~input_layer[1368]),
      .y(Y[510]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron511_1
  function_202 neuron511_1 (
      .a(~input_layer[1338]),
      .b(input_layer[1146]),
      .c(~input_layer[1251]),
      .d(input_layer[1431]),
      .e(input_layer[212]),
      .y(Y[511]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron512_1
  function_26 neuron512_1 (
      .a(input_layer[312]),
      .b(~input_layer[1920]),
      .y(Y[512]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron513_1
  function_40 neuron513_1 (
      .a(~input_layer[1708]),
      .b(~input_layer[975]),
      .c(~input_layer[1026]),
      .d(~input_layer[615]),
      .e(~input_layer[771]),
      .f(~input_layer[512]),
      .y(Y[513]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_203 for neuron514_1
  function_203 neuron514_1 (
      .a(input_layer[2164]),
      .b(~input_layer[384]),
      .c(input_layer[1039]),
      .d(input_layer[614]),
      .e(input_layer[1147]),
      .f(~input_layer[2038]),
      .y(Y[514]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_204 for neuron515_1
  function_204 neuron515_1 (
      .a(~input_layer[1606]),
      .b(~input_layer[460]),
      .c(input_layer[2307]),
      .d(input_layer[1382]),
      .e(~input_layer[1880]),
      .y(Y[515]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron516_1
  function_31 neuron516_1 (
      .a(input_layer[765]),
      .b(input_layer[1436]),
      .c(input_layer[2305]),
      .d(input_layer[938]),
      .e(input_layer[1433]),
      .f(input_layer[670]),
      .y(Y[516]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron517_1
  function_24 neuron517_1 (
      .a(~input_layer[109]),
      .y(Y[517]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron518_1
  function_113 neuron518_1 (
      .a(input_layer[1549]),
      .b(input_layer[2321]),
      .c(input_layer[2287]),
      .d(input_layer[1298]),
      .e(~input_layer[340]),
      .f(~input_layer[1803]),
      .y(Y[518]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron519_1
  function_12 neuron519_1 (
      .a(~input_layer[2087]),
      .b(~input_layer[213]),
      .c(~input_layer[1589]),
      .y(Y[519]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_205 for neuron520_1
  function_205 neuron520_1 (
      .a(input_layer[281]),
      .b(~input_layer[1602]),
      .c(input_layer[1539]),
      .d(~input_layer[1268]),
      .e(~input_layer[1427]),
      .f(input_layer[242]),
      .y(Y[520]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron521_1
  function_14 neuron521_1 (
      .a(~input_layer[998]),
      .b(~input_layer[631]),
      .c(~input_layer[385]),
      .d(~input_layer[984]),
      .e(input_layer[528]),
      .y(Y[521]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_206 for neuron522_1
  function_206 neuron522_1 (
      .a(~input_layer[1914]),
      .b(~input_layer[1318]),
      .c(input_layer[362]),
      .d(input_layer[2215]),
      .e(input_layer[1638]),
      .y(Y[522]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron523_1
  function_44 neuron523_1 (
      .a(~input_layer[1458]),
      .b(input_layer[1189]),
      .c(input_layer[2339]),
      .y(Y[523]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron524_1
  function_132 neuron524_1 (
      .a(input_layer[219]),
      .b(~input_layer[380]),
      .c(~input_layer[889]),
      .d(~input_layer[1404]),
      .e(~input_layer[389]),
      .y(Y[524]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_207 for neuron525_1
  function_207 neuron525_1 (
      .a(~input_layer[1124]),
      .b(input_layer[817]),
      .c(input_layer[940]),
      .d(input_layer[1769]),
      .e(input_layer[809]),
      .f(~input_layer[1526]),
      .y(Y[525]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron526_1
  function_5 neuron526_1 (
      .a(~input_layer[1199]),
      .b(~input_layer[988]),
      .y(Y[526]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron527_1
  function_12 neuron527_1 (
      .a(~input_layer[1572]),
      .b(~input_layer[1003]),
      .c(~input_layer[2166]),
      .y(Y[527]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_208 for neuron528_1
  function_208 neuron528_1 (
      .a(input_layer[1128]),
      .b(~input_layer[2220]),
      .c(~input_layer[1669]),
      .d(~input_layer[1735]),
      .e(input_layer[124]),
      .f(~input_layer[1091]),
      .y(Y[528]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron529_1
  function_63 neuron529_1 (
      .a(input_layer[901]),
      .b(~input_layer[732]),
      .c(input_layer[2166]),
      .d(input_layer[638]),
      .y(Y[529]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_209 for neuron530_1
  function_209 neuron530_1 (
      .a(~input_layer[2153]),
      .b(input_layer[1973]),
      .c(~input_layer[1199]),
      .d(~input_layer[145]),
      .e(input_layer[367]),
      .f(input_layer[1873]),
      .y(Y[530]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron531_1
  function_67 neuron531_1 (
      .a(input_layer[769]),
      .b(~input_layer[985]),
      .c(input_layer[1271]),
      .d(input_layer[1120]),
      .e(~input_layer[1853]),
      .y(Y[531]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron532_1
  function_26 neuron532_1 (
      .a(~input_layer[971]),
      .b(~input_layer[306]),
      .y(Y[532]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron533_1
  function_107 neuron533_1 (
      .a(~input_layer[1053]),
      .b(~input_layer[230]),
      .c(~input_layer[106]),
      .d(~input_layer[1574]),
      .y(Y[533]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron534_1
  function_75 neuron534_1 (
      .a(~input_layer[1618]),
      .b(input_layer[1485]),
      .c(~input_layer[1470]),
      .d(input_layer[2248]),
      .e(~input_layer[1531]),
      .y(Y[534]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron535_1
  function_21 neuron535_1 (
      .a(~input_layer[1469]),
      .b(~input_layer[196]),
      .c(~input_layer[2113]),
      .d(~input_layer[1825]),
      .y(Y[535]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron536_1
  function_67 neuron536_1 (
      .a(input_layer[660]),
      .b(input_layer[1414]),
      .c(~input_layer[2231]),
      .d(input_layer[523]),
      .e(input_layer[1185]),
      .y(Y[536]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron537_1
  function_210 neuron537_1 (
      .a(~input_layer[1668]),
      .b(~input_layer[554]),
      .c(input_layer[232]),
      .d(input_layer[932]),
      .e(input_layer[1689]),
      .y(Y[537]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron538_1
  function_21 neuron538_1 (
      .a(~input_layer[123]),
      .b(input_layer[1393]),
      .c(~input_layer[676]),
      .d(~input_layer[944]),
      .y(Y[538]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron539_1
  function_3 neuron539_1 (
      .a(input_layer[582]),
      .b(input_layer[996]),
      .c(input_layer[1099]),
      .d(input_layer[1539]),
      .e(~input_layer[1558]),
      .y(Y[539]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron540_1
  function_193 neuron540_1 (
      .a(input_layer[270]),
      .b(~input_layer[727]),
      .c(input_layer[973]),
      .d(~input_layer[730]),
      .e(input_layer[622]),
      .f(input_layer[1411]),
      .y(Y[540]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron541_1
  function_148 neuron541_1 (
      .a(~input_layer[195]),
      .b(input_layer[1315]),
      .c(~input_layer[1815]),
      .d(~input_layer[574]),
      .y(Y[541]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron542_1
  function_39 neuron542_1 (
      .a(~input_layer[203]),
      .b(input_layer[648]),
      .c(~input_layer[186]),
      .d(input_layer[534]),
      .y(Y[542]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron543_1
  function_14 neuron543_1 (
      .a(~input_layer[871]),
      .b(~input_layer[136]),
      .c(~input_layer[1639]),
      .d(~input_layer[1512]),
      .e(input_layer[1516]),
      .y(Y[543]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron544_1
  function_3 neuron544_1 (
      .a(input_layer[1445]),
      .b(input_layer[735]),
      .c(input_layer[916]),
      .d(~input_layer[234]),
      .e(input_layer[2058]),
      .y(Y[544]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron545_1
  function_32 neuron545_1 (
      .a(input_layer[1301]),
      .b(~input_layer[377]),
      .c(~input_layer[1246]),
      .d(~input_layer[1880]),
      .y(Y[545]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_143 for neuron546_1
  function_143 neuron546_1 (
      .a(input_layer[612]),
      .b(input_layer[1606]),
      .c(~input_layer[2120]),
      .d(input_layer[909]),
      .e(~input_layer[867]),
      .f(input_layer[1927]),
      .y(Y[546]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_211 for neuron547_1
  function_211 neuron547_1 (
      .a(~input_layer[365]),
      .b(~input_layer[1371]),
      .c(input_layer[2152]),
      .d(~input_layer[1369]),
      .e(~input_layer[673]),
      .y(Y[547]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron548_1
  function_74 neuron548_1 (
      .a(input_layer[379]),
      .b(~input_layer[933]),
      .c(~input_layer[2052]),
      .d(input_layer[780]),
      .e(~input_layer[2338]),
      .y(Y[548]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron549_1
  function_16 neuron549_1 (
      .a(input_layer[1116]),
      .b(input_layer[1409]),
      .c(input_layer[1636]),
      .y(Y[549]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_212 for neuron550_1
  function_212 neuron550_1 (
      .a(input_layer[987]),
      .b(~input_layer[566]),
      .c(input_layer[2067]),
      .d(~input_layer[672]),
      .e(~input_layer[542]),
      .f(input_layer[1858]),
      .y(Y[550]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_213 for neuron551_1
  function_213 neuron551_1 (
      .a(~input_layer[1857]),
      .b(input_layer[2163]),
      .c(~input_layer[1823]),
      .d(~input_layer[1207]),
      .e(input_layer[850]),
      .y(Y[551]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron552_1
  function_26 neuron552_1 (
      .a(input_layer[1555]),
      .b(~input_layer[1711]),
      .y(Y[552]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron553_1
  function_5 neuron553_1 (
      .a(input_layer[484]),
      .b(input_layer[476]),
      .y(Y[553]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron554_1
  function_214 neuron554_1 (
      .a(~input_layer[1438]),
      .b(input_layer[1792]),
      .c(~input_layer[2227]),
      .d(~input_layer[1754]),
      .e(~input_layer[368]),
      .f(input_layer[2046]),
      .y(Y[554]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron555_1
  function_146 neuron555_1 (
      .a(input_layer[2155]),
      .b(input_layer[704]),
      .c(input_layer[442]),
      .d(input_layer[1181]),
      .e(input_layer[1345]),
      .y(Y[555]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron556_1
  function_11 neuron556_1 (
      .a(input_layer[854]),
      .b(input_layer[2089]),
      .c(~input_layer[1032]),
      .d(~input_layer[951]),
      .y(Y[556]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron557_1
  function_53 neuron557_1 (
      .a(input_layer[630]),
      .b(input_layer[1708]),
      .c(~input_layer[1464]),
      .d(~input_layer[1206]),
      .e(~input_layer[1091]),
      .y(Y[557]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_215 for neuron558_1
  function_215 neuron558_1 (
      .a(input_layer[1776]),
      .b(~input_layer[1153]),
      .c(input_layer[1269]),
      .d(input_layer[1961]),
      .e(input_layer[1334]),
      .f(~input_layer[2200]),
      .y(Y[558]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_216 for neuron559_1
  function_216 neuron559_1 (
      .a(input_layer[1281]),
      .b(~input_layer[618]),
      .c(input_layer[311]),
      .d(~input_layer[757]),
      .e(input_layer[567]),
      .f(~input_layer[1426]),
      .y(Y[559]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron560_1
  function_16 neuron560_1 (
      .a(input_layer[394]),
      .b(~input_layer[633]),
      .c(~input_layer[1062]),
      .y(Y[560]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron561_1
  function_45 neuron561_1 (
      .a(~input_layer[1945]),
      .b(input_layer[1132]),
      .c(~input_layer[1947]),
      .d(~input_layer[1641]),
      .e(~input_layer[2074]),
      .f(~input_layer[387]),
      .y(Y[561]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron562_1
  function_20 neuron562_1 (
      .a(input_layer[1199]),
      .b(input_layer[2141]),
      .c(~input_layer[1542]),
      .d(input_layer[348]),
      .e(input_layer[784]),
      .f(input_layer[1847]),
      .y(Y[562]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_217 for neuron563_1
  function_217 neuron563_1 (
      .a(input_layer[1770]),
      .b(~input_layer[1070]),
      .c(~input_layer[1590]),
      .d(~input_layer[399]),
      .e(input_layer[2039]),
      .f(input_layer[1789]),
      .y(Y[563]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[564] = 1'b0;

  // instantiate function_12 for neuron565_1
  function_12 neuron565_1 (
      .a(~input_layer[523]),
      .b(input_layer[1972]),
      .c(~input_layer[1015]),
      .y(Y[565]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron566_1
  function_49 neuron566_1 (
      .a(input_layer[2025]),
      .b(input_layer[1145]),
      .c(input_layer[329]),
      .d(input_layer[670]),
      .e(input_layer[560]),
      .f(input_layer[1563]),
      .y(Y[566]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_218 for neuron567_1
  function_218 neuron567_1 (
      .a(~input_layer[2061]),
      .b(input_layer[300]),
      .c(input_layer[237]),
      .d(input_layer[181]),
      .e(~input_layer[662]),
      .f(~input_layer[987]),
      .y(Y[567]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron568_1
  function_1 neuron568_1 (
      .a(~input_layer[1782]),
      .b(~input_layer[1079]),
      .c(~input_layer[716]),
      .d(input_layer[1040]),
      .e(~input_layer[2169]),
      .f(input_layer[312]),
      .y(Y[568]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron569_1
  function_16 neuron569_1 (
      .a(input_layer[1964]),
      .b(input_layer[904]),
      .c(input_layer[2202]),
      .y(Y[569]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron570_1
  function_76 neuron570_1 (
      .a(~input_layer[1564]),
      .b(~input_layer[779]),
      .c(~input_layer[311]),
      .d(~input_layer[365]),
      .e(~input_layer[459]),
      .f(input_layer[1265]),
      .y(Y[570]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron571_1
  function_10 neuron571_1 (
      .a(input_layer[2135]),
      .b(input_layer[2029]),
      .c(input_layer[1887]),
      .d(~input_layer[1795]),
      .y(Y[571]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron572_1
  function_21 neuron572_1 (
      .a(~input_layer[771]),
      .b(~input_layer[386]),
      .c(~input_layer[1521]),
      .d(~input_layer[1698]),
      .y(Y[572]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron573_1
  function_16 neuron573_1 (
      .a(input_layer[613]),
      .b(input_layer[1916]),
      .c(input_layer[276]),
      .y(Y[573]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_58 for neuron574_1
  function_58 neuron574_1 (
      .a(~input_layer[433]),
      .b(input_layer[549]),
      .c(~input_layer[1561]),
      .d(input_layer[478]),
      .e(input_layer[838]),
      .f(input_layer[828]),
      .y(Y[574]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron575_1
  function_146 neuron575_1 (
      .a(input_layer[2214]),
      .b(~input_layer[1381]),
      .c(input_layer[561]),
      .d(input_layer[885]),
      .e(input_layer[1347]),
      .y(Y[575]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_219 for neuron576_1
  function_219 neuron576_1 (
      .a(~input_layer[2248]),
      .b(input_layer[1254]),
      .c(input_layer[1051]),
      .d(~input_layer[1207]),
      .e(~input_layer[1119]),
      .f(input_layer[1098]),
      .y(Y[576]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron577_1
  function_131 neuron577_1 (
      .a(~input_layer[1872]),
      .b(~input_layer[1877]),
      .c(input_layer[1797]),
      .d(~input_layer[1300]),
      .e(~input_layer[562]),
      .f(~input_layer[545]),
      .y(Y[577]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron578_1
  function_25 neuron578_1 (
      .a(input_layer[985]),
      .b(input_layer[1201]),
      .c(input_layer[787]),
      .d(input_layer[231]),
      .e(input_layer[115]),
      .y(Y[578]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron579_1
  function_16 neuron579_1 (
      .a(input_layer[1374]),
      .b(input_layer[2249]),
      .c(~input_layer[1048]),
      .y(Y[579]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron580_1
  function_42 neuron580_1 (
      .a(input_layer[444]),
      .b(~input_layer[2328]),
      .c(input_layer[2031]),
      .d(~input_layer[99]),
      .e(input_layer[629]),
      .y(Y[580]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron581_1
  function_3 neuron581_1 (
      .a(input_layer[1868]),
      .b(input_layer[2142]),
      .c(input_layer[1187]),
      .d(input_layer[580]),
      .e(input_layer[788]),
      .y(Y[581]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron582_1
  function_5 neuron582_1 (
      .a(input_layer[1183]),
      .b(input_layer[1734]),
      .y(Y[582]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron583_1
  function_63 neuron583_1 (
      .a(input_layer[570]),
      .b(~input_layer[880]),
      .c(input_layer[1157]),
      .d(~input_layer[2315]),
      .y(Y[583]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron584_1
  function_49 neuron584_1 (
      .a(input_layer[1693]),
      .b(input_layer[1949]),
      .c(input_layer[193]),
      .d(~input_layer[1205]),
      .e(~input_layer[981]),
      .f(~input_layer[1594]),
      .y(Y[584]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron585_1
  function_113 neuron585_1 (
      .a(input_layer[2032]),
      .b(input_layer[362]),
      .c(input_layer[323]),
      .d(input_layer[448]),
      .e(input_layer[1333]),
      .f(input_layer[1138]),
      .y(Y[585]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_220 for neuron586_1
  function_220 neuron586_1 (
      .a(input_layer[1956]),
      .b(input_layer[1922]),
      .c(input_layer[1986]),
      .d(input_layer[1978]),
      .e(~input_layer[469]),
      .y(Y[586]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron587_1
  function_221 neuron587_1 (
      .a(~input_layer[2203]),
      .b(~input_layer[1939]),
      .c(~input_layer[634]),
      .d(input_layer[410]),
      .e(~input_layer[411]),
      .f(input_layer[1814]),
      .y(Y[587]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron588_1
  function_17 neuron588_1 (
      .a(~input_layer[1787]),
      .b(~input_layer[825]),
      .c(~input_layer[540]),
      .d(~input_layer[1906]),
      .e(~input_layer[455]),
      .f(~input_layer[34]),
      .y(Y[588]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron589_1
  function_18 neuron589_1 (
      .a(~input_layer[1155]),
      .b(~input_layer[1531]),
      .c(~input_layer[1655]),
      .d(~input_layer[1030]),
      .e(~input_layer[294]),
      .y(Y[589]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_222 for neuron590_1
  function_222 neuron590_1 (
      .a(~input_layer[834]),
      .b(~input_layer[814]),
      .c(~input_layer[2220]),
      .d(~input_layer[660]),
      .e(input_layer[366]),
      .f(input_layer[1815]),
      .y(Y[590]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron591_1
  function_25 neuron591_1 (
      .a(input_layer[1779]),
      .b(input_layer[1135]),
      .c(input_layer[443]),
      .d(input_layer[1649]),
      .e(input_layer[1860]),
      .y(Y[591]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron592_1
  function_169 neuron592_1 (
      .a(input_layer[1052]),
      .b(input_layer[2025]),
      .c(input_layer[1473]),
      .d(input_layer[774]),
      .e(~input_layer[399]),
      .f(~input_layer[365]),
      .y(Y[592]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_223 for neuron593_1
  function_223 neuron593_1 (
      .a(~input_layer[760]),
      .b(input_layer[1729]),
      .c(~input_layer[2230]),
      .d(input_layer[328]),
      .e(input_layer[1645]),
      .f(input_layer[1717]),
      .y(Y[593]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron594_1
  function_32 neuron594_1 (
      .a(input_layer[1466]),
      .b(input_layer[1130]),
      .c(~input_layer[2330]),
      .d(~input_layer[1043]),
      .y(Y[594]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron595_1
  function_12 neuron595_1 (
      .a(~input_layer[1586]),
      .b(~input_layer[454]),
      .c(~input_layer[1909]),
      .y(Y[595]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron596_1
  function_221 neuron596_1 (
      .a(~input_layer[1370]),
      .b(~input_layer[1308]),
      .c(~input_layer[1400]),
      .d(input_layer[1815]),
      .e(~input_layer[940]),
      .f(input_layer[2054]),
      .y(Y[596]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron597_1
  function_12 neuron597_1 (
      .a(~input_layer[1128]),
      .b(~input_layer[2200]),
      .c(~input_layer[2225]),
      .y(Y[597]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron598_1
  function_53 neuron598_1 (
      .a(input_layer[455]),
      .b(input_layer[1916]),
      .c(input_layer[566]),
      .d(~input_layer[2304]),
      .e(~input_layer[1392]),
      .y(Y[598]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_224 for neuron599_1
  function_224 neuron599_1 (
      .a(~input_layer[1373]),
      .b(~input_layer[1211]),
      .c(input_layer[775]),
      .d(input_layer[711]),
      .y(Y[599]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_225 for neuron600_1
  function_225 neuron600_1 (
      .a(~input_layer[1546]),
      .b(input_layer[1819]),
      .c(input_layer[1938]),
      .d(~input_layer[202]),
      .e(input_layer[1846]),
      .f(input_layer[1007]),
      .y(Y[600]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron601_1
  function_20 neuron601_1 (
      .a(input_layer[1672]),
      .b(input_layer[2290]),
      .c(~input_layer[450]),
      .d(input_layer[1593]),
      .e(~input_layer[2032]),
      .f(input_layer[1802]),
      .y(Y[601]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron602_1
  function_4 neuron602_1 (
      .a(input_layer[388]),
      .b(input_layer[1762]),
      .c(~input_layer[2193]),
      .d(input_layer[1807]),
      .e(input_layer[2011]),
      .y(Y[602]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron603_1
  function_93 neuron603_1 (
      .a(~input_layer[1337]),
      .b(~input_layer[2157]),
      .c(input_layer[884]),
      .d(~input_layer[469]),
      .e(~input_layer[2291]),
      .f(input_layer[1715]),
      .y(Y[603]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_195 for neuron604_1
  function_195 neuron604_1 (
      .a(input_layer[395]),
      .b(input_layer[1667]),
      .c(~input_layer[731]),
      .d(~input_layer[2319]),
      .e(input_layer[2254]),
      .f(input_layer[1432]),
      .y(Y[604]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron605_1
  function_3 neuron605_1 (
      .a(input_layer[301]),
      .b(input_layer[1274]),
      .c(input_layer[2146]),
      .d(~input_layer[1899]),
      .e(input_layer[1396]),
      .y(Y[605]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron606_1
  function_16 neuron606_1 (
      .a(input_layer[197]),
      .b(input_layer[865]),
      .c(input_layer[2076]),
      .y(Y[606]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron607_1
  function_135 neuron607_1 (
      .a(~input_layer[2139]),
      .b(input_layer[1889]),
      .c(input_layer[1448]),
      .d(~input_layer[1311]),
      .e(input_layer[1994]),
      .y(Y[607]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_42 for neuron608_1
  function_42 neuron608_1 (
      .a(~input_layer[300]),
      .b(input_layer[2166]),
      .c(input_layer[1691]),
      .d(input_layer[1517]),
      .e(~input_layer[1906]),
      .y(Y[608]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron609_1
  function_21 neuron609_1 (
      .a(~input_layer[298]),
      .b(input_layer[1290]),
      .c(~input_layer[1674]),
      .d(~input_layer[1856]),
      .y(Y[609]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron610_1
  function_49 neuron610_1 (
      .a(input_layer[2118]),
      .b(input_layer[1837]),
      .c(input_layer[1017]),
      .d(~input_layer[962]),
      .e(input_layer[1103]),
      .f(input_layer[1852]),
      .y(Y[610]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron611_1
  function_67 neuron611_1 (
      .a(input_layer[2039]),
      .b(input_layer[123]),
      .c(input_layer[109]),
      .d(~input_layer[1556]),
      .e(~input_layer[996]),
      .y(Y[611]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron612_1
  function_3 neuron612_1 (
      .a(input_layer[1368]),
      .b(input_layer[1836]),
      .c(input_layer[764]),
      .d(~input_layer[607]),
      .e(~input_layer[1617]),
      .y(Y[612]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_8 for neuron613_1
  function_8 neuron613_1 (
      .a(~input_layer[1052]),
      .b(~input_layer[271]),
      .c(input_layer[640]),
      .d(~input_layer[1746]),
      .e(~input_layer[467]),
      .f(input_layer[1177]),
      .y(Y[613]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron614_1
  function_76 neuron614_1 (
      .a(~input_layer[474]),
      .b(~input_layer[658]),
      .c(~input_layer[1526]),
      .d(~input_layer[1863]),
      .e(~input_layer[1549]),
      .f(~input_layer[1971]),
      .y(Y[614]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron615_1
  function_99 neuron615_1 (
      .a(input_layer[1647]),
      .b(input_layer[1537]),
      .c(input_layer[1581]),
      .d(input_layer[936]),
      .e(input_layer[1237]),
      .f(input_layer[1943]),
      .y(Y[615]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron616_1
  function_152 neuron616_1 (
      .a(~input_layer[686]),
      .b(input_layer[638]),
      .c(input_layer[806]),
      .d(~input_layer[2308]),
      .e(input_layer[1492]),
      .f(~input_layer[1301]),
      .y(Y[616]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron617_1
  function_107 neuron617_1 (
      .a(~input_layer[625]),
      .b(~input_layer[437]),
      .c(~input_layer[1603]),
      .d(input_layer[2198]),
      .y(Y[617]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron618_1
  function_18 neuron618_1 (
      .a(~input_layer[1890]),
      .b(~input_layer[1504]),
      .c(~input_layer[598]),
      .d(~input_layer[850]),
      .e(~input_layer[1448]),
      .y(Y[618]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_226 for neuron619_1
  function_226 neuron619_1 (
      .a(~input_layer[1582]),
      .b(input_layer[2207]),
      .c(input_layer[787]),
      .d(~input_layer[439]),
      .e(input_layer[149]),
      .f(~input_layer[436]),
      .y(Y[619]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_227 for neuron620_1
  function_227 neuron620_1 (
      .a(~input_layer[579]),
      .b(input_layer[1120]),
      .c(~input_layer[669]),
      .d(input_layer[1217]),
      .e(~input_layer[695]),
      .f(input_layer[1679]),
      .y(Y[620]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_228 for neuron621_1
  function_228 neuron621_1 (
      .a(~input_layer[1700]),
      .b(input_layer[218]),
      .c(input_layer[116]),
      .d(~input_layer[784]),
      .e(~input_layer[1084]),
      .f(input_layer[134]),
      .y(Y[621]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_229 for neuron622_1
  function_229 neuron622_1 (
      .a(~input_layer[911]),
      .b(input_layer[596]),
      .c(input_layer[1264]),
      .d(~input_layer[1893]),
      .e(~input_layer[1698]),
      .f(input_layer[331]),
      .y(Y[622]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_230 for neuron623_1
  function_230 neuron623_1 (
      .a(~input_layer[1470]),
      .b(~input_layer[2167]),
      .c(input_layer[701]),
      .d(~input_layer[1503]),
      .e(input_layer[1206]),
      .f(~input_layer[664]),
      .y(Y[623]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron624_1
  function_231 neuron624_1 (
      .a(input_layer[552]),
      .b(~input_layer[1915]),
      .c(input_layer[908]),
      .d(~input_layer[2178]),
      .e(~input_layer[1021]),
      .f(~input_layer[1958]),
      .y(Y[624]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron625_1
  function_3 neuron625_1 (
      .a(input_layer[472]),
      .b(input_layer[1279]),
      .c(input_layer[2003]),
      .d(~input_layer[846]),
      .e(~input_layer[1555]),
      .y(Y[625]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron626_1
  function_232 neuron626_1 (
      .a(~input_layer[1045]),
      .b(input_layer[1146]),
      .c(input_layer[887]),
      .d(input_layer[763]),
      .e(~input_layer[1829]),
      .y(Y[626]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron627_1
  function_92 neuron627_1 (
      .a(~input_layer[491]),
      .b(~input_layer[1207]),
      .c(input_layer[184]),
      .d(input_layer[2125]),
      .y(Y[627]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron628_1
  function_148 neuron628_1 (
      .a(~input_layer[2129]),
      .b(input_layer[1722]),
      .c(input_layer[469]),
      .d(~input_layer[2256]),
      .y(Y[628]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_233 for neuron629_1
  function_233 neuron629_1 (
      .a(~input_layer[1624]),
      .b(input_layer[2051]),
      .c(~input_layer[2314]),
      .d(~input_layer[1486]),
      .e(~input_layer[1322]),
      .f(~input_layer[504]),
      .y(Y[629]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron630_1
  function_234 neuron630_1 (
      .a(~input_layer[1587]),
      .b(~input_layer[788]),
      .c(~input_layer[2005]),
      .d(input_layer[520]),
      .e(input_layer[1804]),
      .f(~input_layer[831]),
      .y(Y[630]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron631_1
  function_49 neuron631_1 (
      .a(input_layer[1871]),
      .b(input_layer[2241]),
      .c(input_layer[2230]),
      .d(input_layer[2161]),
      .e(input_layer[1813]),
      .f(input_layer[814]),
      .y(Y[631]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron632_1
  function_202 neuron632_1 (
      .a(~input_layer[1203]),
      .b(input_layer[883]),
      .c(input_layer[769]),
      .d(~input_layer[532]),
      .e(input_layer[551]),
      .y(Y[632]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron633_1
  function_32 neuron633_1 (
      .a(~input_layer[987]),
      .b(input_layer[301]),
      .c(~input_layer[949]),
      .d(~input_layer[1608]),
      .y(Y[633]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron634_1
  function_18 neuron634_1 (
      .a(~input_layer[1834]),
      .b(~input_layer[1326]),
      .c(~input_layer[1463]),
      .d(~input_layer[123]),
      .e(~input_layer[1685]),
      .y(Y[634]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_160 for neuron635_1
  function_160 neuron635_1 (
      .a(input_layer[323]),
      .b(input_layer[1387]),
      .c(~input_layer[724]),
      .d(input_layer[1461]),
      .e(~input_layer[990]),
      .y(Y[635]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_213 for neuron636_1
  function_213 neuron636_1 (
      .a(~input_layer[115]),
      .b(input_layer[539]),
      .c(~input_layer[113]),
      .d(~input_layer[1122]),
      .e(input_layer[537]),
      .y(Y[636]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron637_1
  function_169 neuron637_1 (
      .a(input_layer[1158]),
      .b(input_layer[1422]),
      .c(input_layer[1301]),
      .d(input_layer[426]),
      .e(~input_layer[732]),
      .f(~input_layer[2257]),
      .y(Y[637]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron638_1
  function_11 neuron638_1 (
      .a(input_layer[1154]),
      .b(input_layer[2251]),
      .c(input_layer[1599]),
      .d(input_layer[1094]),
      .y(Y[638]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron639_1
  function_18 neuron639_1 (
      .a(~input_layer[1726]),
      .b(~input_layer[599]),
      .c(~input_layer[514]),
      .d(~input_layer[1853]),
      .e(input_layer[723]),
      .y(Y[639]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron640_1
  function_92 neuron640_1 (
      .a(~input_layer[1200]),
      .b(input_layer[1254]),
      .c(input_layer[604]),
      .d(~input_layer[112]),
      .y(Y[640]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron641_1
  function_48 neuron641_1 (
      .a(input_layer[2046]),
      .b(input_layer[2083]),
      .c(~input_layer[1490]),
      .d(input_layer[482]),
      .e(input_layer[1515]),
      .y(Y[641]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron642_1
  function_149 neuron642_1 (
      .a(~input_layer[1082]),
      .b(~input_layer[949]),
      .c(~input_layer[865]),
      .d(~input_layer[837]),
      .y(Y[642]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron643_1
  function_18 neuron643_1 (
      .a(~input_layer[832]),
      .b(~input_layer[679]),
      .c(~input_layer[1083]),
      .d(~input_layer[1810]),
      .e(~input_layer[345]),
      .y(Y[643]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron644_1
  function_67 neuron644_1 (
      .a(input_layer[724]),
      .b(input_layer[1960]),
      .c(input_layer[889]),
      .d(~input_layer[1657]),
      .e(~input_layer[990]),
      .y(Y[644]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron645_1
  function_44 neuron645_1 (
      .a(input_layer[303]),
      .b(~input_layer[2074]),
      .c(~input_layer[1231]),
      .y(Y[645]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron646_1
  function_21 neuron646_1 (
      .a(~input_layer[718]),
      .b(~input_layer[1016]),
      .c(~input_layer[669]),
      .d(input_layer[1116]),
      .y(Y[646]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron647_1
  function_11 neuron647_1 (
      .a(input_layer[1244]),
      .b(input_layer[2119]),
      .c(input_layer[1775]),
      .d(~input_layer[889]),
      .y(Y[647]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron648_1
  function_18 neuron648_1 (
      .a(~input_layer[1058]),
      .b(~input_layer[464]),
      .c(~input_layer[276]),
      .d(~input_layer[1744]),
      .e(~input_layer[1941]),
      .y(Y[648]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron649_1
  function_35 neuron649_1 (
      .a(~input_layer[1978]),
      .b(~input_layer[1688]),
      .c(input_layer[2202]),
      .d(~input_layer[502]),
      .e(~input_layer[41]),
      .y(Y[649]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron650_1
  function_92 neuron650_1 (
      .a(input_layer[405]),
      .b(~input_layer[1893]),
      .c(~input_layer[1330]),
      .d(~input_layer[877]),
      .y(Y[650]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron651_1
  function_112 neuron651_1 (
      .a(~input_layer[472]),
      .b(~input_layer[440]),
      .c(input_layer[1018]),
      .d(input_layer[804]),
      .e(~input_layer[1408]),
      .f(input_layer[1359]),
      .y(Y[651]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron652_1
  function_53 neuron652_1 (
      .a(input_layer[2035]),
      .b(input_layer[883]),
      .c(input_layer[2286]),
      .d(input_layer[1899]),
      .e(input_layer[1361]),
      .y(Y[652]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron653_1
  function_12 neuron653_1 (
      .a(~input_layer[1075]),
      .b(~input_layer[368]),
      .c(~input_layer[1083]),
      .y(Y[653]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron654_1
  function_12 neuron654_1 (
      .a(~input_layer[1231]),
      .b(~input_layer[230]),
      .c(input_layer[1323]),
      .y(Y[654]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron655_1
  function_18 neuron655_1 (
      .a(~input_layer[1022]),
      .b(~input_layer[1256]),
      .c(input_layer[878]),
      .d(~input_layer[1754]),
      .e(~input_layer[262]),
      .y(Y[655]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron656_1
  function_120 neuron656_1 (
      .a(~input_layer[714]),
      .b(~input_layer[1153]),
      .c(input_layer[741]),
      .d(input_layer[1121]),
      .e(~input_layer[1913]),
      .f(~input_layer[1101]),
      .y(Y[656]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_235 for neuron657_1
  function_235 neuron657_1 (
      .a(~input_layer[1381]),
      .b(~input_layer[359]),
      .c(~input_layer[1371]),
      .d(input_layer[2330]),
      .e(input_layer[2147]),
      .f(~input_layer[1596]),
      .y(Y[657]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron658_1
  function_21 neuron658_1 (
      .a(~input_layer[952]),
      .b(~input_layer[214]),
      .c(input_layer[543]),
      .d(~input_layer[2245]),
      .y(Y[658]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron659_1
  function_31 neuron659_1 (
      .a(input_layer[1698]),
      .b(input_layer[1733]),
      .c(input_layer[769]),
      .d(input_layer[1899]),
      .e(input_layer[1996]),
      .f(input_layer[1915]),
      .y(Y[659]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_215 for neuron660_1
  function_215 neuron660_1 (
      .a(input_layer[2160]),
      .b(~input_layer[1778]),
      .c(~input_layer[1816]),
      .d(input_layer[1290]),
      .e(input_layer[2175]),
      .f(~input_layer[1296]),
      .y(Y[660]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron661_1
  function_193 neuron661_1 (
      .a(input_layer[1994]),
      .b(input_layer[2318]),
      .c(~input_layer[803]),
      .d(~input_layer[1530]),
      .e(~input_layer[553]),
      .f(input_layer[1325]),
      .y(Y[661]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron662_1
  function_63 neuron662_1 (
      .a(input_layer[1132]),
      .b(~input_layer[1039]),
      .c(input_layer[1568]),
      .d(input_layer[152]),
      .y(Y[662]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron663_1
  function_148 neuron663_1 (
      .a(~input_layer[1744]),
      .b(input_layer[881]),
      .c(~input_layer[1066]),
      .d(input_layer[1117]),
      .y(Y[663]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron664_1
  function_179 neuron664_1 (
      .a(~input_layer[1190]),
      .b(input_layer[271]),
      .c(~input_layer[1360]),
      .d(input_layer[962]),
      .e(input_layer[405]),
      .y(Y[664]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron665_1
  function_26 neuron665_1 (
      .a(~input_layer[2154]),
      .b(~input_layer[1616]),
      .y(Y[665]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_236 for neuron666_1
  function_236 neuron666_1 (
      .a(~input_layer[1106]),
      .b(input_layer[288]),
      .c(input_layer[468]),
      .d(input_layer[1547]),
      .e(~input_layer[2247]),
      .f(~input_layer[1849]),
      .y(Y[666]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron667_1
  function_95 neuron667_1 (
      .a(input_layer[2287]),
      .b(input_layer[1737]),
      .c(input_layer[797]),
      .d(~input_layer[1913]),
      .y(Y[667]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron668_1
  function_44 neuron668_1 (
      .a(~input_layer[1491]),
      .b(input_layer[702]),
      .c(input_layer[1573]),
      .y(Y[668]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron669_1
  function_0 neuron669_1 (
      .a(input_layer[1362]),
      .b(input_layer[1755]),
      .c(input_layer[1454]),
      .d(~input_layer[837]),
      .e(input_layer[448]),
      .y(Y[669]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_237 for neuron670_1
  function_237 neuron670_1 (
      .a(input_layer[483]),
      .b(~input_layer[2231]),
      .c(~input_layer[893]),
      .d(input_layer[241]),
      .e(input_layer[99]),
      .f(input_layer[545]),
      .y(Y[670]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron671_1
  function_76 neuron671_1 (
      .a(~input_layer[381]),
      .b(~input_layer[446]),
      .c(~input_layer[1943]),
      .d(~input_layer[2027]),
      .e(input_layer[553]),
      .f(~input_layer[2283]),
      .y(Y[671]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron672_1
  function_0 neuron672_1 (
      .a(~input_layer[1969]),
      .b(input_layer[1016]),
      .c(input_layer[1271]),
      .d(input_layer[306]),
      .e(input_layer[957]),
      .y(Y[672]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_238 for neuron673_1
  function_238 neuron673_1 (
      .a(input_layer[1885]),
      .b(~input_layer[496]),
      .c(~input_layer[1258]),
      .d(~input_layer[969]),
      .e(input_layer[1028]),
      .y(Y[673]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron674_1
  function_95 neuron674_1 (
      .a(~input_layer[1554]),
      .b(input_layer[991]),
      .c(input_layer[961]),
      .d(~input_layer[1843]),
      .y(Y[674]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron675_1
  function_116 neuron675_1 (
      .a(input_layer[679]),
      .b(input_layer[1844]),
      .c(input_layer[730]),
      .d(~input_layer[452]),
      .y(Y[675]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron676_1
  function_10 neuron676_1 (
      .a(input_layer[1482]),
      .b(input_layer[537]),
      .c(~input_layer[1018]),
      .d(input_layer[1537]),
      .y(Y[676]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron677_1
  function_91 neuron677_1 (
      .a(input_layer[1613]),
      .b(input_layer[203]),
      .c(~input_layer[704]),
      .d(input_layer[1769]),
      .e(input_layer[2077]),
      .f(~input_layer[758]),
      .y(Y[677]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_239 for neuron678_1
  function_239 neuron678_1 (
      .a(input_layer[1656]),
      .b(input_layer[267]),
      .c(input_layer[2254]),
      .d(~input_layer[404]),
      .e(~input_layer[1147]),
      .y(Y[678]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_240 for neuron679_1
  function_240 neuron679_1 (
      .a(input_layer[728]),
      .b(~input_layer[920]),
      .c(input_layer[432]),
      .d(input_layer[1877]),
      .e(~input_layer[669]),
      .f(~input_layer[1778]),
      .y(Y[679]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron680_1
  function_241 neuron680_1 (
      .a(~input_layer[2042]),
      .b(input_layer[1386]),
      .c(input_layer[904]),
      .d(input_layer[851]),
      .e(input_layer[1120]),
      .f(~input_layer[773]),
      .y(Y[680]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron681_1
  function_63 neuron681_1 (
      .a(input_layer[2203]),
      .b(~input_layer[1079]),
      .c(~input_layer[1966]),
      .d(~input_layer[1540]),
      .y(Y[681]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron682_1
  function_11 neuron682_1 (
      .a(input_layer[2141]),
      .b(input_layer[1084]),
      .c(~input_layer[1460]),
      .d(input_layer[718]),
      .y(Y[682]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron683_1
  function_26 neuron683_1 (
      .a(~input_layer[1666]),
      .b(~input_layer[469]),
      .y(Y[683]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron684_1
  function_16 neuron684_1 (
      .a(input_layer[737]),
      .b(input_layer[2073]),
      .c(input_layer[1675]),
      .y(Y[684]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_109 for neuron685_1
  function_109 neuron685_1 (
      .a(input_layer[1547]),
      .b(input_layer[1218]),
      .c(input_layer[293]),
      .d(~input_layer[2296]),
      .e(input_layer[120]),
      .f(input_layer[2228]),
      .y(Y[685]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron686_1
  function_234 neuron686_1 (
      .a(~input_layer[1612]),
      .b(~input_layer[1923]),
      .c(~input_layer[1908]),
      .d(~input_layer[660]),
      .e(input_layer[2171]),
      .f(input_layer[543]),
      .y(Y[686]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron687_1
  function_149 neuron687_1 (
      .a(~input_layer[2230]),
      .b(~input_layer[1606]),
      .c(input_layer[993]),
      .d(input_layer[1111]),
      .y(Y[687]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron688_1
  function_95 neuron688_1 (
      .a(input_layer[2035]),
      .b(input_layer[2134]),
      .c(~input_layer[1989]),
      .d(~input_layer[153]),
      .y(Y[688]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron689_1
  function_113 neuron689_1 (
      .a(~input_layer[1966]),
      .b(input_layer[296]),
      .c(input_layer[286]),
      .d(input_layer[1475]),
      .e(input_layer[1149]),
      .f(input_layer[1257]),
      .y(Y[689]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_242 for neuron690_1
  function_242 neuron690_1 (
      .a(input_layer[872]),
      .b(~input_layer[1867]),
      .c(~input_layer[374]),
      .d(~input_layer[324]),
      .e(input_layer[905]),
      .f(input_layer[1237]),
      .y(Y[690]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron691_1
  function_24 neuron691_1 (
      .a(input_layer[1961]),
      .y(Y[691]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron692_1
  function_32 neuron692_1 (
      .a(input_layer[1209]),
      .b(~input_layer[2198]),
      .c(input_layer[405]),
      .d(input_layer[1037]),
      .y(Y[692]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron693_1
  function_113 neuron693_1 (
      .a(input_layer[662]),
      .b(input_layer[830]),
      .c(input_layer[1083]),
      .d(input_layer[1549]),
      .e(input_layer[713]),
      .f(input_layer[1982]),
      .y(Y[693]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron694_1
  function_92 neuron694_1 (
      .a(input_layer[2006]),
      .b(~input_layer[977]),
      .c(~input_layer[1604]),
      .d(input_layer[815]),
      .y(Y[694]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_112 for neuron695_1
  function_112 neuron695_1 (
      .a(~input_layer[1412]),
      .b(~input_layer[1902]),
      .c(~input_layer[1012]),
      .d(input_layer[1520]),
      .e(~input_layer[1942]),
      .f(~input_layer[843]),
      .y(Y[695]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[696] = 1'b0;

  // instantiate function_10 for neuron697_1
  function_10 neuron697_1 (
      .a(input_layer[1783]),
      .b(input_layer[433]),
      .c(input_layer[659]),
      .d(input_layer[909]),
      .y(Y[697]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_243 for neuron698_1
  function_243 neuron698_1 (
      .a(input_layer[1163]),
      .b(~input_layer[619]),
      .c(~input_layer[1059]),
      .d(~input_layer[1003]),
      .e(input_layer[1606]),
      .f(input_layer[1414]),
      .y(Y[698]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron699_1
  function_113 neuron699_1 (
      .a(input_layer[574]),
      .b(input_layer[646]),
      .c(input_layer[2233]),
      .d(~input_layer[308]),
      .e(~input_layer[1546]),
      .f(input_layer[1172]),
      .y(Y[699]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron700_1
  function_148 neuron700_1 (
      .a(~input_layer[1299]),
      .b(~input_layer[1416]),
      .c(~input_layer[2156]),
      .d(input_layer[785]),
      .y(Y[700]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron701_1
  function_14 neuron701_1 (
      .a(~input_layer[1127]),
      .b(~input_layer[1282]),
      .c(~input_layer[2166]),
      .d(input_layer[2123]),
      .e(~input_layer[1645]),
      .y(Y[701]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_244 for neuron702_1
  function_244 neuron702_1 (
      .a(input_layer[193]),
      .b(~input_layer[2003]),
      .c(input_layer[1096]),
      .d(~input_layer[1035]),
      .e(input_layer[729]),
      .f(input_layer[2338]),
      .y(Y[702]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron703_1
  function_107 neuron703_1 (
      .a(input_layer[904]),
      .b(~input_layer[754]),
      .c(~input_layer[886]),
      .d(input_layer[473]),
      .y(Y[703]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron704_1
  function_3 neuron704_1 (
      .a(input_layer[850]),
      .b(input_layer[1588]),
      .c(input_layer[2160]),
      .d(~input_layer[886]),
      .e(input_layer[722]),
      .y(Y[704]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_245 for neuron705_1
  function_245 neuron705_1 (
      .a(input_layer[1549]),
      .b(~input_layer[1907]),
      .c(~input_layer[1644]),
      .d(input_layer[1719]),
      .e(input_layer[2032]),
      .f(input_layer[1768]),
      .y(Y[705]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron706_1
  function_16 neuron706_1 (
      .a(input_layer[2206]),
      .b(~input_layer[1146]),
      .c(~input_layer[1395]),
      .y(Y[706]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron707_1
  function_67 neuron707_1 (
      .a(input_layer[1244]),
      .b(input_layer[975]),
      .c(~input_layer[951]),
      .d(input_layer[2326]),
      .e(input_layer[2096]),
      .y(Y[707]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron708_1
  function_10 neuron708_1 (
      .a(input_layer[1801]),
      .b(input_layer[713]),
      .c(~input_layer[609]),
      .d(input_layer[2089]),
      .y(Y[708]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron709_1
  function_167 neuron709_1 (
      .a(~input_layer[288]),
      .b(input_layer[859]),
      .c(~input_layer[380]),
      .d(input_layer[1278]),
      .e(input_layer[1478]),
      .y(Y[709]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron710_1
  function_11 neuron710_1 (
      .a(input_layer[1664]),
      .b(input_layer[309]),
      .c(input_layer[2218]),
      .d(input_layer[234]),
      .y(Y[710]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_55 for neuron711_1
  function_55 neuron711_1 (
      .a(~input_layer[1647]),
      .b(~input_layer[752]),
      .c(input_layer[717]),
      .d(input_layer[1113]),
      .e(input_layer[271]),
      .f(~input_layer[1295]),
      .y(Y[711]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron712_1
  function_18 neuron712_1 (
      .a(~input_layer[206]),
      .b(~input_layer[1816]),
      .c(~input_layer[2296]),
      .d(~input_layer[1939]),
      .e(~input_layer[1604]),
      .y(Y[712]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_246 for neuron713_1
  function_246 neuron713_1 (
      .a(input_layer[1610]),
      .b(~input_layer[2314]),
      .c(input_layer[1947]),
      .d(~input_layer[1126]),
      .e(~input_layer[412]),
      .f(~input_layer[654]),
      .y(Y[713]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron714_1
  function_95 neuron714_1 (
      .a(~input_layer[1049]),
      .b(input_layer[1336]),
      .c(input_layer[1328]),
      .d(~input_layer[1571]),
      .y(Y[714]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron715_1
  function_14 neuron715_1 (
      .a(~input_layer[451]),
      .b(input_layer[1149]),
      .c(~input_layer[675]),
      .d(~input_layer[1600]),
      .e(~input_layer[1509]),
      .y(Y[715]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_247 for neuron716_1
  function_247 neuron716_1 (
      .a(~input_layer[664]),
      .b(~input_layer[1801]),
      .c(input_layer[2049]),
      .d(~input_layer[1443]),
      .e(input_layer[2335]),
      .y(Y[716]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron717_1
  function_76 neuron717_1 (
      .a(~input_layer[1717]),
      .b(~input_layer[201]),
      .c(~input_layer[195]),
      .d(~input_layer[2236]),
      .e(input_layer[1602]),
      .f(~input_layer[1940]),
      .y(Y[717]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron718_1
  function_248 neuron718_1 (
      .a(~input_layer[2249]),
      .b(input_layer[1470]),
      .c(~input_layer[2319]),
      .d(~input_layer[2202]),
      .e(~input_layer[648]),
      .f(input_layer[893]),
      .y(Y[718]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_249 for neuron719_1
  function_249 neuron719_1 (
      .a(~input_layer[1906]),
      .b(input_layer[2214]),
      .c(input_layer[1578]),
      .d(input_layer[2322]),
      .e(input_layer[1185]),
      .f(~input_layer[1602]),
      .y(Y[719]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron720_1
  function_12 neuron720_1 (
      .a(~input_layer[1673]),
      .b(~input_layer[1357]),
      .c(input_layer[958]),
      .y(Y[720]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron721_1
  function_113 neuron721_1 (
      .a(input_layer[627]),
      .b(input_layer[2142]),
      .c(~input_layer[1140]),
      .d(input_layer[929]),
      .e(input_layer[717]),
      .f(~input_layer[1764]),
      .y(Y[721]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron722_1
  function_5 neuron722_1 (
      .a(input_layer[1543]),
      .b(input_layer[2318]),
      .y(Y[722]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron723_1
  function_24 neuron723_1 (
      .a(~input_layer[1303]),
      .y(Y[723]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron724_1
  function_74 neuron724_1 (
      .a(input_layer[1972]),
      .b(~input_layer[1288]),
      .c(~input_layer[1820]),
      .d(input_layer[890]),
      .e(input_layer[987]),
      .y(Y[724]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_250 for neuron725_1
  function_250 neuron725_1 (
      .a(input_layer[1588]),
      .b(input_layer[299]),
      .c(input_layer[444]),
      .d(~input_layer[2337]),
      .e(input_layer[1770]),
      .f(input_layer[1439]),
      .y(Y[725]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron726_1
  function_11 neuron726_1 (
      .a(input_layer[1799]),
      .b(input_layer[226]),
      .c(~input_layer[1219]),
      .d(input_layer[1416]),
      .y(Y[726]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_251 for neuron727_1
  function_251 neuron727_1 (
      .a(input_layer[324]),
      .b(input_layer[1892]),
      .c(~input_layer[1385]),
      .d(~input_layer[525]),
      .e(input_layer[2280]),
      .f(input_layer[327]),
      .y(Y[727]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron728_1
  function_10 neuron728_1 (
      .a(input_layer[448]),
      .b(input_layer[1567]),
      .c(input_layer[1733]),
      .d(input_layer[1158]),
      .y(Y[728]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_252 for neuron729_1
  function_252 neuron729_1 (
      .a(~input_layer[207]),
      .b(input_layer[1014]),
      .c(input_layer[1247]),
      .d(input_layer[518]),
      .e(input_layer[1952]),
      .f(~input_layer[2234]),
      .y(Y[729]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_222 for neuron730_1
  function_222 neuron730_1 (
      .a(input_layer[991]),
      .b(input_layer[1112]),
      .c(~input_layer[1314]),
      .d(~input_layer[1838]),
      .e(input_layer[1616]),
      .f(input_layer[728]),
      .y(Y[730]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron731_1
  function_253 neuron731_1 (
      .a(~input_layer[485]),
      .b(input_layer[734]),
      .c(input_layer[775]),
      .d(input_layer[2336]),
      .e(input_layer[2072]),
      .y(Y[731]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_254 for neuron732_1
  function_254 neuron732_1 (
      .a(~input_layer[1786]),
      .b(~input_layer[1658]),
      .c(input_layer[885]),
      .d(~input_layer[1710]),
      .e(~input_layer[1304]),
      .f(input_layer[852]),
      .y(Y[732]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron733_1
  function_100 neuron733_1 (
      .a(input_layer[556]),
      .b(input_layer[1831]),
      .c(~input_layer[1984]),
      .y(Y[733]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron734_1
  function_1 neuron734_1 (
      .a(~input_layer[1400]),
      .b(~input_layer[217]),
      .c(~input_layer[2011]),
      .d(input_layer[702]),
      .e(~input_layer[1513]),
      .f(input_layer[2098]),
      .y(Y[734]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_255 for neuron735_1
  function_255 neuron735_1 (
      .a(input_layer[2234]),
      .b(input_layer[2117]),
      .c(input_layer[2333]),
      .d(~input_layer[1666]),
      .e(~input_layer[1150]),
      .y(Y[735]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron736_1
  function_61 neuron736_1 (
      .a(~input_layer[1548]),
      .b(input_layer[1882]),
      .c(input_layer[1966]),
      .d(input_layer[2155]),
      .e(~input_layer[486]),
      .y(Y[736]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_220 for neuron737_1
  function_220 neuron737_1 (
      .a(input_layer[513]),
      .b(input_layer[2122]),
      .c(~input_layer[298]),
      .d(input_layer[1108]),
      .e(~input_layer[1128]),
      .y(Y[737]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron738_1
  function_45 neuron738_1 (
      .a(~input_layer[867]),
      .b(~input_layer[1435]),
      .c(~input_layer[1103]),
      .d(~input_layer[1940]),
      .e(~input_layer[379]),
      .f(~input_layer[1708]),
      .y(Y[738]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron739_1
  function_107 neuron739_1 (
      .a(~input_layer[1789]),
      .b(~input_layer[1489]),
      .c(~input_layer[731]),
      .d(~input_layer[601]),
      .y(Y[739]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron740_1
  function_34 neuron740_1 (
      .a(input_layer[296]),
      .b(~input_layer[1396]),
      .c(~input_layer[1022]),
      .d(input_layer[1853]),
      .e(input_layer[1157]),
      .y(Y[740]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron741_1
  function_44 neuron741_1 (
      .a(~input_layer[767]),
      .b(input_layer[1050]),
      .c(~input_layer[1198]),
      .y(Y[741]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron742_1
  function_14 neuron742_1 (
      .a(~input_layer[968]),
      .b(~input_layer[410]),
      .c(~input_layer[1079]),
      .d(input_layer[1701]),
      .e(input_layer[1780]),
      .y(Y[742]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron743_1
  function_18 neuron743_1 (
      .a(~input_layer[1503]),
      .b(~input_layer[1229]),
      .c(~input_layer[1568]),
      .d(~input_layer[911]),
      .e(~input_layer[1983]),
      .y(Y[743]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron744_1
  function_125 neuron744_1 (
      .a(~input_layer[2319]),
      .b(input_layer[954]),
      .c(input_layer[903]),
      .d(~input_layer[1348]),
      .e(~input_layer[1976]),
      .y(Y[744]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_6 for neuron745_1
  function_6 neuron745_1 (
      .a(~input_layer[919]),
      .b(input_layer[2239]),
      .c(~input_layer[1040]),
      .d(input_layer[327]),
      .e(input_layer[1928]),
      .f(input_layer[1485]),
      .y(Y[745]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron746_1
  function_34 neuron746_1 (
      .a(input_layer[651]),
      .b(input_layer[1983]),
      .c(~input_layer[1549]),
      .d(input_layer[972]),
      .e(~input_layer[479]),
      .y(Y[746]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_73 for neuron747_1
  function_73 neuron747_1 (
      .a(~input_layer[999]),
      .b(input_layer[225]),
      .c(input_layer[2317]),
      .d(input_layer[979]),
      .e(~input_layer[1818]),
      .f(input_layer[1316]),
      .y(Y[747]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron748_1
  function_24 neuron748_1 (
      .a(input_layer[811]),
      .y(Y[748]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron749_1
  function_10 neuron749_1 (
      .a(input_layer[431]),
      .b(~input_layer[1459]),
      .c(~input_layer[1624]),
      .d(~input_layer[1865]),
      .y(Y[749]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_256 for neuron750_1
  function_256 neuron750_1 (
      .a(input_layer[1974]),
      .b(input_layer[111]),
      .c(~input_layer[302]),
      .d(~input_layer[2096]),
      .e(input_layer[1773]),
      .y(Y[750]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron751_1
  function_25 neuron751_1 (
      .a(input_layer[1775]),
      .b(input_layer[2125]),
      .c(input_layer[853]),
      .d(input_layer[959]),
      .e(input_layer[1603]),
      .y(Y[751]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron752_1
  function_16 neuron752_1 (
      .a(input_layer[990]),
      .b(input_layer[1320]),
      .c(input_layer[2036]),
      .y(Y[752]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_257 for neuron753_1
  function_257 neuron753_1 (
      .a(input_layer[767]),
      .b(~input_layer[1732]),
      .c(~input_layer[517]),
      .d(input_layer[694]),
      .e(~input_layer[240]),
      .y(Y[753]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron754_1
  function_100 neuron754_1 (
      .a(input_layer[2165]),
      .b(input_layer[558]),
      .c(input_layer[634]),
      .y(Y[754]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_258 for neuron755_1
  function_258 neuron755_1 (
      .a(input_layer[811]),
      .b(~input_layer[200]),
      .c(~input_layer[1628]),
      .d(input_layer[884]),
      .e(input_layer[1004]),
      .f(~input_layer[1323]),
      .y(Y[755]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron756_1
  function_12 neuron756_1 (
      .a(~input_layer[899]),
      .b(~input_layer[1697]),
      .c(input_layer[482]),
      .y(Y[756]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_59 for neuron757_1
  function_59 neuron757_1 (
      .a(~input_layer[486]),
      .b(~input_layer[1783]),
      .c(input_layer[2286]),
      .d(input_layer[806]),
      .e(input_layer[642]),
      .f(input_layer[1554]),
      .y(Y[757]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron758_1
  function_30 neuron758_1 (
      .a(~input_layer[1065]),
      .b(input_layer[1745]),
      .c(input_layer[1645]),
      .d(input_layer[1426]),
      .y(Y[758]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron759_1
  function_61 neuron759_1 (
      .a(input_layer[1216]),
      .b(~input_layer[1534]),
      .c(input_layer[1668]),
      .d(~input_layer[560]),
      .e(input_layer[2113]),
      .y(Y[759]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron760_1
  function_149 neuron760_1 (
      .a(~input_layer[688]),
      .b(input_layer[752]),
      .c(~input_layer[1767]),
      .d(~input_layer[122]),
      .y(Y[760]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_237 for neuron761_1
  function_237 neuron761_1 (
      .a(~input_layer[1340]),
      .b(input_layer[2223]),
      .c(~input_layer[1695]),
      .d(input_layer[2289]),
      .e(input_layer[1273]),
      .f(~input_layer[374]),
      .y(Y[761]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_259 for neuron762_1
  function_259 neuron762_1 (
      .a(input_layer[1047]),
      .b(input_layer[1506]),
      .c(~input_layer[565]),
      .d(~input_layer[503]),
      .e(~input_layer[618]),
      .f(~input_layer[2186]),
      .y(Y[762]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron763_1
  function_63 neuron763_1 (
      .a(~input_layer[1381]),
      .b(input_layer[2310]),
      .c(~input_layer[1902]),
      .d(~input_layer[1154]),
      .y(Y[763]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron764_1
  function_49 neuron764_1 (
      .a(input_layer[1234]),
      .b(input_layer[1571]),
      .c(input_layer[684]),
      .d(input_layer[1151]),
      .e(input_layer[120]),
      .f(input_layer[1947]),
      .y(Y[764]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron765_1
  function_61 neuron765_1 (
      .a(~input_layer[903]),
      .b(input_layer[551]),
      .c(~input_layer[777]),
      .d(~input_layer[593]),
      .e(~input_layer[1745]),
      .y(Y[765]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron766_1
  function_11 neuron766_1 (
      .a(input_layer[318]),
      .b(input_layer[1327]),
      .c(input_layer[2245]),
      .d(input_layer[1230]),
      .y(Y[766]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron767_1
  function_67 neuron767_1 (
      .a(input_layer[1157]),
      .b(input_layer[2007]),
      .c(input_layer[187]),
      .d(input_layer[2169]),
      .e(~input_layer[728]),
      .y(Y[767]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron768_1
  function_116 neuron768_1 (
      .a(input_layer[1779]),
      .b(input_layer[1657]),
      .c(input_layer[1410]),
      .d(input_layer[522]),
      .y(Y[768]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron769_1
  function_24 neuron769_1 (
      .a(~input_layer[1962]),
      .y(Y[769]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron770_1
  function_107 neuron770_1 (
      .a(~input_layer[1566]),
      .b(~input_layer[1642]),
      .c(~input_layer[838]),
      .d(input_layer[2336]),
      .y(Y[770]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_260 for neuron771_1
  function_260 neuron771_1 (
      .a(input_layer[1464]),
      .b(~input_layer[888]),
      .c(~input_layer[1854]),
      .d(~input_layer[1137]),
      .e(input_layer[1140]),
      .f(input_layer[38]),
      .y(Y[771]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[772] = 1'b0;

  // instantiate function_154 for neuron773_1
  function_154 neuron773_1 (
      .a(input_layer[2147]),
      .b(input_layer[1468]),
      .c(input_layer[1231]),
      .d(input_layer[776]),
      .e(~input_layer[1203]),
      .y(Y[773]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron774_1
  function_167 neuron774_1 (
      .a(~input_layer[1991]),
      .b(input_layer[614]),
      .c(input_layer[1572]),
      .d(~input_layer[635]),
      .e(input_layer[1363]),
      .y(Y[774]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron775_1
  function_44 neuron775_1 (
      .a(~input_layer[1217]),
      .b(~input_layer[302]),
      .c(input_layer[2290]),
      .y(Y[775]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron776_1
  function_11 neuron776_1 (
      .a(input_layer[1754]),
      .b(input_layer[792]),
      .c(~input_layer[1891]),
      .d(input_layer[918]),
      .y(Y[776]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron777_1
  function_64 neuron777_1 (
      .a(input_layer[718]),
      .b(input_layer[2306]),
      .c(~input_layer[863]),
      .d(input_layer[309]),
      .e(input_layer[1106]),
      .y(Y[777]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron778_1
  function_56 neuron778_1 (
      .a(~input_layer[1632]),
      .b(~input_layer[1606]),
      .c(input_layer[1239]),
      .d(input_layer[793]),
      .e(~input_layer[2200]),
      .y(Y[778]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_70 for neuron779_1
  function_70 neuron779_1 (
      .a(input_layer[1741]),
      .b(~input_layer[845]),
      .c(~input_layer[484]),
      .d(~input_layer[430]),
      .e(~input_layer[1392]),
      .f(~input_layer[273]),
      .y(Y[779]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_261 for neuron780_1
  function_261 neuron780_1 (
      .a(~input_layer[1650]),
      .b(input_layer[1392]),
      .c(~input_layer[2035]),
      .d(input_layer[1205]),
      .e(~input_layer[368]),
      .f(input_layer[1756]),
      .y(Y[780]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron781_1
  function_12 neuron781_1 (
      .a(~input_layer[1116]),
      .b(~input_layer[1842]),
      .c(~input_layer[1721]),
      .y(Y[781]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron782_1
  function_232 neuron782_1 (
      .a(~input_layer[2306]),
      .b(input_layer[2215]),
      .c(input_layer[238]),
      .d(input_layer[1773]),
      .e(input_layer[1922]),
      .y(Y[782]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron783_1
  function_33 neuron783_1 (
      .a(~input_layer[599]),
      .b(~input_layer[1505]),
      .c(~input_layer[1590]),
      .d(input_layer[2052]),
      .e(input_layer[625]),
      .y(Y[783]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron784_1
  function_89 neuron784_1 (
      .a(~input_layer[2134]),
      .b(input_layer[128]),
      .c(input_layer[1184]),
      .d(input_layer[139]),
      .e(~input_layer[1035]),
      .f(~input_layer[1455]),
      .y(Y[784]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_262 for neuron785_1
  function_262 neuron785_1 (
      .a(input_layer[1589]),
      .b(input_layer[395]),
      .c(~input_layer[1894]),
      .d(input_layer[1026]),
      .e(~input_layer[1534]),
      .f(input_layer[578]),
      .y(Y[785]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron786_1
  function_92 neuron786_1 (
      .a(input_layer[543]),
      .b(~input_layer[718]),
      .c(~input_layer[759]),
      .d(~input_layer[514]),
      .y(Y[786]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron787_1
  function_10 neuron787_1 (
      .a(input_layer[1472]),
      .b(input_layer[2161]),
      .c(input_layer[593]),
      .d(~input_layer[1893]),
      .y(Y[787]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron788_1
  function_0 neuron788_1 (
      .a(input_layer[600]),
      .b(input_layer[1253]),
      .c(input_layer[1145]),
      .d(input_layer[1481]),
      .e(~input_layer[956]),
      .y(Y[788]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron789_1
  function_170 neuron789_1 (
      .a(~input_layer[641]),
      .b(~input_layer[1250]),
      .c(input_layer[2167]),
      .d(input_layer[1640]),
      .e(~input_layer[123]),
      .y(Y[789]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron790_1
  function_17 neuron790_1 (
      .a(~input_layer[1589]),
      .b(~input_layer[1172]),
      .c(input_layer[2251]),
      .d(input_layer[735]),
      .e(~input_layer[1565]),
      .f(~input_layer[11]),
      .y(Y[790]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron791_1
  function_172 neuron791_1 (
      .a(~input_layer[460]),
      .b(input_layer[2202]),
      .c(~input_layer[2166]),
      .d(input_layer[2130]),
      .e(input_layer[706]),
      .f(~input_layer[794]),
      .y(Y[791]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron792_1
  function_21 neuron792_1 (
      .a(~input_layer[2060]),
      .b(~input_layer[2306]),
      .c(~input_layer[615]),
      .d(~input_layer[2150]),
      .y(Y[792]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron793_1
  function_175 neuron793_1 (
      .a(~input_layer[640]),
      .b(input_layer[2313]),
      .c(~input_layer[122]),
      .d(input_layer[1302]),
      .e(~input_layer[607]),
      .y(Y[793]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron794_1
  function_148 neuron794_1 (
      .a(~input_layer[405]),
      .b(input_layer[803]),
      .c(input_layer[598]),
      .d(~input_layer[981]),
      .y(Y[794]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron795_1
  function_5 neuron795_1 (
      .a(~input_layer[1363]),
      .b(input_layer[969]),
      .y(Y[795]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron796_1
  function_19 neuron796_1 (
      .a(~input_layer[1969]),
      .b(input_layer[1147]),
      .c(input_layer[2076]),
      .d(~input_layer[895]),
      .y(Y[796]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron797_1
  function_18 neuron797_1 (
      .a(~input_layer[1580]),
      .b(~input_layer[1405]),
      .c(~input_layer[516]),
      .d(~input_layer[763]),
      .e(~input_layer[1267]),
      .y(Y[797]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_263 for neuron798_1
  function_263 neuron798_1 (
      .a(~input_layer[1912]),
      .b(~input_layer[1206]),
      .c(input_layer[2304]),
      .d(~input_layer[1976]),
      .e(input_layer[928]),
      .f(input_layer[601]),
      .y(Y[798]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron799_1
  function_37 neuron799_1 (
      .a(input_layer[306]),
      .b(~input_layer[1320]),
      .c(input_layer[1492]),
      .d(input_layer[1341]),
      .e(input_layer[2011]),
      .y(Y[799]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron800_1
  function_11 neuron800_1 (
      .a(input_layer[1355]),
      .b(input_layer[2208]),
      .c(input_layer[2116]),
      .d(input_layer[348]),
      .y(Y[800]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron801_1
  function_25 neuron801_1 (
      .a(input_layer[481]),
      .b(input_layer[556]),
      .c(input_layer[1753]),
      .d(input_layer[680]),
      .e(input_layer[525]),
      .y(Y[801]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_264 for neuron802_1
  function_264 neuron802_1 (
      .a(~input_layer[560]),
      .b(~input_layer[1943]),
      .c(input_layer[127]),
      .d(input_layer[1168]),
      .e(input_layer[195]),
      .f(input_layer[130]),
      .y(Y[802]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron803_1
  function_56 neuron803_1 (
      .a(~input_layer[1126]),
      .b(~input_layer[1739]),
      .c(~input_layer[1243]),
      .d(~input_layer[103]),
      .e(~input_layer[1610]),
      .y(Y[803]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron804_1
  function_107 neuron804_1 (
      .a(~input_layer[581]),
      .b(input_layer[636]),
      .c(~input_layer[1493]),
      .d(input_layer[855]),
      .y(Y[804]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron805_1
  function_25 neuron805_1 (
      .a(input_layer[1365]),
      .b(input_layer[1909]),
      .c(input_layer[1868]),
      .d(~input_layer[1274]),
      .e(~input_layer[1315]),
      .y(Y[805]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron806_1
  function_11 neuron806_1 (
      .a(input_layer[2223]),
      .b(input_layer[770]),
      .c(input_layer[144]),
      .d(~input_layer[1396]),
      .y(Y[806]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron807_1
  function_91 neuron807_1 (
      .a(input_layer[632]),
      .b(input_layer[238]),
      .c(~input_layer[569]),
      .d(input_layer[2085]),
      .e(~input_layer[947]),
      .f(input_layer[1461]),
      .y(Y[807]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron808_1
  function_130 neuron808_1 (
      .a(~input_layer[1113]),
      .b(~input_layer[1447]),
      .c(input_layer[511]),
      .d(input_layer[1929]),
      .e(~input_layer[350]),
      .f(~input_layer[170]),
      .y(Y[808]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron809_1
  function_119 neuron809_1 (
      .a(input_layer[1112]),
      .b(input_layer[139]),
      .c(input_layer[2144]),
      .d(~input_layer[1447]),
      .e(~input_layer[1670]),
      .f(input_layer[1610]),
      .y(Y[809]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron810_1
  function_25 neuron810_1 (
      .a(input_layer[1660]),
      .b(input_layer[1697]),
      .c(input_layer[2146]),
      .d(input_layer[599]),
      .e(input_layer[731]),
      .y(Y[810]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron811_1
  function_10 neuron811_1 (
      .a(input_layer[1300]),
      .b(input_layer[2317]),
      .c(input_layer[325]),
      .d(~input_layer[720]),
      .y(Y[811]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_220 for neuron812_1
  function_220 neuron812_1 (
      .a(input_layer[1549]),
      .b(input_layer[1463]),
      .c(input_layer[1115]),
      .d(input_layer[1001]),
      .e(~input_layer[1770]),
      .y(Y[812]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_85 for neuron813_1
  function_85 neuron813_1 (
      .a(input_layer[298]),
      .b(~input_layer[348]),
      .c(input_layer[141]),
      .d(input_layer[860]),
      .e(~input_layer[1571]),
      .f(input_layer[816]),
      .y(Y[813]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron814_1
  function_40 neuron814_1 (
      .a(~input_layer[802]),
      .b(~input_layer[767]),
      .c(input_layer[474]),
      .d(~input_layer[515]),
      .e(~input_layer[1683]),
      .f(~input_layer[1440]),
      .y(Y[814]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_265 for neuron815_1
  function_265 neuron815_1 (
      .a(input_layer[1459]),
      .b(input_layer[239]),
      .c(~input_layer[845]),
      .d(~input_layer[1182]),
      .e(~input_layer[1011]),
      .f(input_layer[2107]),
      .y(Y[815]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron816_1
  function_104 neuron816_1 (
      .a(input_layer[2208]),
      .b(~input_layer[574]),
      .c(~input_layer[1034]),
      .y(Y[816]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron817_1
  function_3 neuron817_1 (
      .a(input_layer[2124]),
      .b(input_layer[115]),
      .c(input_layer[838]),
      .d(input_layer[1318]),
      .e(input_layer[2241]),
      .y(Y[817]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron818_1
  function_44 neuron818_1 (
      .a(~input_layer[1363]),
      .b(input_layer[1217]),
      .c(~input_layer[2079]),
      .y(Y[818]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron819_1
  function_146 neuron819_1 (
      .a(input_layer[1703]),
      .b(input_layer[538]),
      .c(~input_layer[1296]),
      .d(~input_layer[1222]),
      .e(~input_layer[960]),
      .y(Y[819]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_98 for neuron820_1
  function_98 neuron820_1 (
      .a(input_layer[2026]),
      .b(~input_layer[617]),
      .c(input_layer[191]),
      .d(~input_layer[1288]),
      .e(~input_layer[275]),
      .y(Y[820]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[821] = 1'b1;

  // instantiate function_139 for neuron822_1
  function_139 neuron822_1 (
      .a(input_layer[1607]),
      .b(~input_layer[568]),
      .c(input_layer[884]),
      .d(input_layer[261]),
      .e(input_layer[1892]),
      .y(Y[822]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron823_1
  function_16 neuron823_1 (
      .a(~input_layer[727]),
      .b(input_layer[495]),
      .c(input_layer[2023]),
      .y(Y[823]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_266 for neuron824_1
  function_266 neuron824_1 (
      .a(~input_layer[741]),
      .b(~input_layer[2328]),
      .c(input_layer[1522]),
      .d(~input_layer[128]),
      .e(input_layer[693]),
      .f(input_layer[18]),
      .y(Y[824]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron825_1
  function_100 neuron825_1 (
      .a(input_layer[2141]),
      .b(~input_layer[1800]),
      .c(input_layer[702]),
      .y(Y[825]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron826_1
  function_12 neuron826_1 (
      .a(~input_layer[916]),
      .b(~input_layer[880]),
      .c(~input_layer[232]),
      .y(Y[826]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_267 for neuron827_1
  function_267 neuron827_1 (
      .a(~input_layer[1629]),
      .b(input_layer[104]),
      .c(input_layer[473]),
      .d(input_layer[798]),
      .e(~input_layer[203]),
      .f(~input_layer[1698]),
      .y(Y[827]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_268 for neuron828_1
  function_268 neuron828_1 (
      .a(~input_layer[2249]),
      .b(~input_layer[1057]),
      .c(~input_layer[883]),
      .d(input_layer[1819]),
      .e(~input_layer[1982]),
      .f(input_layer[70]),
      .y(Y[828]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron829_1
  function_167 neuron829_1 (
      .a(~input_layer[572]),
      .b(input_layer[2134]),
      .c(input_layer[282]),
      .d(input_layer[1238]),
      .e(~input_layer[1176]),
      .y(Y[829]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron830_1
  function_132 neuron830_1 (
      .a(~input_layer[386]),
      .b(input_layer[218]),
      .c(input_layer[1100]),
      .d(input_layer[897]),
      .e(~input_layer[545]),
      .y(Y[830]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron831_1
  function_148 neuron831_1 (
      .a(input_layer[1120]),
      .b(~input_layer[143]),
      .c(input_layer[1230]),
      .d(input_layer[385]),
      .y(Y[831]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_269 for neuron832_1
  function_269 neuron832_1 (
      .a(input_layer[2086]),
      .b(~input_layer[697]),
      .c(~input_layer[1084]),
      .d(~input_layer[887]),
      .e(~input_layer[1258]),
      .f(input_layer[227]),
      .y(Y[832]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron833_1
  function_32 neuron833_1 (
      .a(input_layer[1711]),
      .b(~input_layer[1533]),
      .c(input_layer[240]),
      .d(input_layer[1491]),
      .y(Y[833]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_270 for neuron834_1
  function_270 neuron834_1 (
      .a(input_layer[1965]),
      .b(input_layer[2032]),
      .c(input_layer[453]),
      .d(~input_layer[1208]),
      .e(~input_layer[2073]),
      .f(~input_layer[2257]),
      .y(Y[834]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron835_1
  function_61 neuron835_1 (
      .a(~input_layer[692]),
      .b(input_layer[1373]),
      .c(input_layer[1728]),
      .d(~input_layer[986]),
      .e(input_layer[1800]),
      .y(Y[835]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron836_1
  function_44 neuron836_1 (
      .a(~input_layer[537]),
      .b(~input_layer[1056]),
      .c(~input_layer[351]),
      .y(Y[836]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron837_1
  function_61 neuron837_1 (
      .a(~input_layer[200]),
      .b(input_layer[1124]),
      .c(~input_layer[1632]),
      .d(input_layer[1644]),
      .e(input_layer[1538]),
      .y(Y[837]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron838_1
  function_67 neuron838_1 (
      .a(input_layer[1732]),
      .b(input_layer[1488]),
      .c(input_layer[1149]),
      .d(~input_layer[1473]),
      .e(input_layer[2093]),
      .y(Y[838]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron839_1
  function_17 neuron839_1 (
      .a(~input_layer[628]),
      .b(~input_layer[1777]),
      .c(~input_layer[1275]),
      .d(input_layer[1332]),
      .e(~input_layer[348]),
      .f(~input_layer[2038]),
      .y(Y[839]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron840_1
  function_37 neuron840_1 (
      .a(input_layer[1161]),
      .b(~input_layer[658]),
      .c(input_layer[682]),
      .d(input_layer[105]),
      .e(input_layer[316]),
      .y(Y[840]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron841_1
  function_26 neuron841_1 (
      .a(~input_layer[308]),
      .b(~input_layer[1011]),
      .y(Y[841]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron842_1
  function_12 neuron842_1 (
      .a(~input_layer[1358]),
      .b(~input_layer[1199]),
      .c(input_layer[1537]),
      .y(Y[842]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_271 for neuron843_1
  function_271 neuron843_1 (
      .a(input_layer[791]),
      .b(~input_layer[199]),
      .c(input_layer[2205]),
      .d(~input_layer[2251]),
      .e(~input_layer[1089]),
      .f(~input_layer[260]),
      .y(Y[843]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron844_1
  function_21 neuron844_1 (
      .a(~input_layer[1146]),
      .b(~input_layer[1487]),
      .c(~input_layer[851]),
      .d(~input_layer[2319]),
      .y(Y[844]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_208 for neuron845_1
  function_208 neuron845_1 (
      .a(~input_layer[1716]),
      .b(~input_layer[272]),
      .c(input_layer[1874]),
      .d(~input_layer[2317]),
      .e(~input_layer[134]),
      .f(~input_layer[263]),
      .y(Y[845]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_272 for neuron846_1
  function_272 neuron846_1 (
      .a(input_layer[1278]),
      .b(~input_layer[1137]),
      .c(~input_layer[842]),
      .d(~input_layer[1406]),
      .e(input_layer[982]),
      .f(input_layer[167]),
      .y(Y[846]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron847_1
  function_107 neuron847_1 (
      .a(~input_layer[1970]),
      .b(~input_layer[950]),
      .c(input_layer[102]),
      .d(~input_layer[1433]),
      .y(Y[847]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron848_1
  function_21 neuron848_1 (
      .a(~input_layer[1590]),
      .b(~input_layer[193]),
      .c(~input_layer[1363]),
      .d(input_layer[1047]),
      .y(Y[848]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron849_1
  function_90 neuron849_1 (
      .a(~input_layer[720]),
      .b(~input_layer[1686]),
      .c(input_layer[607]),
      .d(~input_layer[261]),
      .e(input_layer[2081]),
      .y(Y[849]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron850_1
  function_139 neuron850_1 (
      .a(~input_layer[966]),
      .b(input_layer[2196]),
      .c(input_layer[798]),
      .d(input_layer[330]),
      .e(input_layer[2096]),
      .y(Y[850]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron851_1
  function_130 neuron851_1 (
      .a(input_layer[785]),
      .b(input_layer[1080]),
      .c(~input_layer[1985]),
      .d(input_layer[1765]),
      .e(input_layer[339]),
      .f(input_layer[58]),
      .y(Y[851]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron852_1
  function_11 neuron852_1 (
      .a(input_layer[297]),
      .b(input_layer[436]),
      .c(input_layer[1749]),
      .d(input_layer[596]),
      .y(Y[852]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_262 for neuron853_1
  function_262 neuron853_1 (
      .a(input_layer[220]),
      .b(~input_layer[1107]),
      .c(input_layer[1672]),
      .d(input_layer[2338]),
      .e(~input_layer[2085]),
      .f(~input_layer[338]),
      .y(Y[853]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron854_1
  function_11 neuron854_1 (
      .a(input_layer[599]),
      .b(input_layer[935]),
      .c(input_layer[1252]),
      .d(~input_layer[2149]),
      .y(Y[854]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron855_1
  function_21 neuron855_1 (
      .a(~input_layer[2168]),
      .b(~input_layer[128]),
      .c(input_layer[871]),
      .d(input_layer[1736]),
      .y(Y[855]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron856_1
  function_16 neuron856_1 (
      .a(input_layer[2134]),
      .b(input_layer[1814]),
      .c(input_layer[219]),
      .y(Y[856]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_273 for neuron857_1
  function_273 neuron857_1 (
      .a(~input_layer[147]),
      .b(input_layer[2117]),
      .c(~input_layer[1538]),
      .d(~input_layer[1075]),
      .e(~input_layer[1736]),
      .f(input_layer[841]),
      .y(Y[857]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron858_1
  function_11 neuron858_1 (
      .a(input_layer[206]),
      .b(input_layer[1021]),
      .c(input_layer[716]),
      .d(input_layer[2173]),
      .y(Y[858]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_274 for neuron859_1
  function_274 neuron859_1 (
      .a(input_layer[2304]),
      .b(~input_layer[402]),
      .c(~input_layer[955]),
      .d(~input_layer[1990]),
      .e(~input_layer[873]),
      .f(input_layer[1847]),
      .y(Y[859]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_247 for neuron860_1
  function_247 neuron860_1 (
      .a(~input_layer[209]),
      .b(input_layer[2060]),
      .c(~input_layer[1202]),
      .d(~input_layer[1482]),
      .e(~input_layer[1401]),
      .y(Y[860]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_275 for neuron861_1
  function_275 neuron861_1 (
      .a(input_layer[965]),
      .b(input_layer[1041]),
      .c(~input_layer[1831]),
      .d(~input_layer[1187]),
      .e(input_layer[1214]),
      .f(~input_layer[1873]),
      .y(Y[861]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron862_1
  function_44 neuron862_1 (
      .a(input_layer[1360]),
      .b(~input_layer[2214]),
      .c(input_layer[2122]),
      .y(Y[862]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron863_1
  function_24 neuron863_1 (
      .a(input_layer[1059]),
      .y(Y[863]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_276 for neuron864_1
  function_276 neuron864_1 (
      .a(input_layer[950]),
      .b(~input_layer[548]),
      .c(~input_layer[2203]),
      .d(~input_layer[2246]),
      .e(~input_layer[100]),
      .y(Y[864]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron865_1
  function_16 neuron865_1 (
      .a(input_layer[870]),
      .b(~input_layer[1957]),
      .c(input_layer[2114]),
      .y(Y[865]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_277 for neuron866_1
  function_277 neuron866_1 (
      .a(~input_layer[988]),
      .b(input_layer[597]),
      .c(~input_layer[1602]),
      .d(input_layer[1758]),
      .e(~input_layer[1294]),
      .y(Y[866]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron867_1
  function_146 neuron867_1 (
      .a(input_layer[1473]),
      .b(input_layer[1354]),
      .c(~input_layer[863]),
      .d(input_layer[2111]),
      .e(~input_layer[839]),
      .y(Y[867]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron868_1
  function_31 neuron868_1 (
      .a(input_layer[911]),
      .b(input_layer[600]),
      .c(input_layer[1777]),
      .d(input_layer[586]),
      .e(input_layer[2334]),
      .f(input_layer[2043]),
      .y(Y[868]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_131 for neuron869_1
  function_131 neuron869_1 (
      .a(~input_layer[1390]),
      .b(input_layer[1141]),
      .c(~input_layer[794]),
      .d(~input_layer[595]),
      .e(input_layer[2022]),
      .f(~input_layer[378]),
      .y(Y[869]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron870_1
  function_107 neuron870_1 (
      .a(~input_layer[1745]),
      .b(input_layer[1041]),
      .c(~input_layer[118]),
      .d(input_layer[1240]),
      .y(Y[870]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron871_1
  function_49 neuron871_1 (
      .a(input_layer[776]),
      .b(input_layer[1482]),
      .c(input_layer[837]),
      .d(input_layer[197]),
      .e(input_layer[982]),
      .f(input_layer[2283]),
      .y(Y[871]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron872_1
  function_76 neuron872_1 (
      .a(~input_layer[1135]),
      .b(~input_layer[1755]),
      .c(~input_layer[1295]),
      .d(~input_layer[1909]),
      .e(~input_layer[428]),
      .f(~input_layer[1222]),
      .y(Y[872]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron873_1
  function_139 neuron873_1 (
      .a(input_layer[1506]),
      .b(input_layer[1396]),
      .c(~input_layer[2301]),
      .d(input_layer[2194]),
      .e(~input_layer[642]),
      .y(Y[873]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron874_1
  function_125 neuron874_1 (
      .a(~input_layer[2034]),
      .b(~input_layer[2326]),
      .c(~input_layer[1924]),
      .d(input_layer[1939]),
      .e(~input_layer[1845]),
      .y(Y[874]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron875_1
  function_107 neuron875_1 (
      .a(~input_layer[993]),
      .b(~input_layer[764]),
      .c(~input_layer[2155]),
      .d(input_layer[645]),
      .y(Y[875]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron876_1
  function_162 neuron876_1 (
      .a(~input_layer[1864]),
      .b(~input_layer[712]),
      .c(input_layer[1410]),
      .d(~input_layer[1443]),
      .e(~input_layer[1854]),
      .y(Y[876]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron877_1
  function_24 neuron877_1 (
      .a(~input_layer[1893]),
      .y(Y[877]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron878_1
  function_35 neuron878_1 (
      .a(~input_layer[214]),
      .b(~input_layer[1570]),
      .c(~input_layer[1217]),
      .d(input_layer[1748]),
      .e(~input_layer[1649]),
      .y(Y[878]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron879_1
  function_170 neuron879_1 (
      .a(~input_layer[1587]),
      .b(input_layer[1101]),
      .c(~input_layer[548]),
      .d(~input_layer[1425]),
      .e(input_layer[2143]),
      .y(Y[879]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_278 for neuron880_1
  function_278 neuron880_1 (
      .a(input_layer[1902]),
      .b(~input_layer[692]),
      .c(input_layer[1453]),
      .d(input_layer[638]),
      .e(~input_layer[2243]),
      .f(~input_layer[620]),
      .y(Y[880]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_279 for neuron881_1
  function_279 neuron881_1 (
      .a(~input_layer[482]),
      .b(input_layer[2227]),
      .c(~input_layer[405]),
      .d(input_layer[1591]),
      .e(input_layer[1350]),
      .y(Y[881]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_36 for neuron882_1
  function_36 neuron882_1 (
      .a(~input_layer[2318]),
      .b(input_layer[1363]),
      .c(input_layer[1725]),
      .d(~input_layer[2326]),
      .e(input_layer[180]),
      .f(input_layer[1006]),
      .y(Y[882]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron883_1
  function_17 neuron883_1 (
      .a(~input_layer[2125]),
      .b(~input_layer[284]),
      .c(input_layer[962]),
      .d(~input_layer[1470]),
      .e(input_layer[912]),
      .f(input_layer[535]),
      .y(Y[883]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_244 for neuron884_1
  function_244 neuron884_1 (
      .a(~input_layer[822]),
      .b(input_layer[1841]),
      .c(input_layer[106]),
      .d(input_layer[397]),
      .e(input_layer[579]),
      .f(~input_layer[946]),
      .y(Y[884]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron885_1
  function_10 neuron885_1 (
      .a(~input_layer[1150]),
      .b(~input_layer[1384]),
      .c(input_layer[934]),
      .d(~input_layer[1724]),
      .y(Y[885]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron886_1
  function_130 neuron886_1 (
      .a(input_layer[1030]),
      .b(input_layer[1075]),
      .c(input_layer[1545]),
      .d(~input_layer[1663]),
      .e(~input_layer[739]),
      .f(input_layer[318]),
      .y(Y[886]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_280 for neuron887_1
  function_280 neuron887_1 (
      .a(input_layer[940]),
      .b(input_layer[2227]),
      .c(~input_layer[464]),
      .d(input_layer[2112]),
      .e(input_layer[1519]),
      .f(~input_layer[46]),
      .y(Y[887]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_281 for neuron888_1
  function_281 neuron888_1 (
      .a(input_layer[1359]),
      .b(~input_layer[1424]),
      .c(~input_layer[1558]),
      .d(~input_layer[1914]),
      .e(input_layer[1099]),
      .f(~input_layer[689]),
      .y(Y[888]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron889_1
  function_202 neuron889_1 (
      .a(input_layer[995]),
      .b(~input_layer[216]),
      .c(~input_layer[1126]),
      .d(~input_layer[868]),
      .e(~input_layer[1313]),
      .y(Y[889]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron890_1
  function_11 neuron890_1 (
      .a(input_layer[1620]),
      .b(input_layer[696]),
      .c(input_layer[142]),
      .d(~input_layer[1307]),
      .y(Y[890]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_282 for neuron891_1
  function_282 neuron891_1 (
      .a(~input_layer[131]),
      .b(input_layer[814]),
      .c(input_layer[818]),
      .d(~input_layer[1622]),
      .e(input_layer[184]),
      .y(Y[891]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron892_1
  function_53 neuron892_1 (
      .a(input_layer[721]),
      .b(input_layer[843]),
      .c(input_layer[717]),
      .d(input_layer[2250]),
      .e(~input_layer[1390]),
      .y(Y[892]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron893_1
  function_12 neuron893_1 (
      .a(~input_layer[1449]),
      .b(~input_layer[2247]),
      .c(~input_layer[1639]),
      .y(Y[893]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron894_1
  function_21 neuron894_1 (
      .a(~input_layer[1395]),
      .b(~input_layer[777]),
      .c(~input_layer[2305]),
      .d(~input_layer[1351]),
      .y(Y[894]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron895_1
  function_113 neuron895_1 (
      .a(input_layer[1353]),
      .b(~input_layer[1117]),
      .c(input_layer[1001]),
      .d(input_layer[296]),
      .e(input_layer[732]),
      .f(input_layer[502]),
      .y(Y[895]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_88 for neuron896_1
  function_88 neuron896_1 (
      .a(~input_layer[1193]),
      .b(input_layer[1583]),
      .c(input_layer[353]),
      .d(input_layer[532]),
      .e(input_layer[483]),
      .f(~input_layer[141]),
      .y(Y[896]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron897_1
  function_10 neuron897_1 (
      .a(input_layer[1779]),
      .b(input_layer[931]),
      .c(~input_layer[823]),
      .d(~input_layer[563]),
      .y(Y[897]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_283 for neuron898_1
  function_283 neuron898_1 (
      .a(input_layer[1951]),
      .b(~input_layer[986]),
      .c(~input_layer[1087]),
      .d(input_layer[1984]),
      .e(~input_layer[2344]),
      .f(~input_layer[82]),
      .y(Y[898]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron899_1
  function_44 neuron899_1 (
      .a(~input_layer[870]),
      .b(~input_layer[1164]),
      .c(~input_layer[1531]),
      .y(Y[899]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron900_1
  function_154 neuron900_1 (
      .a(input_layer[847]),
      .b(input_layer[1634]),
      .c(~input_layer[2080]),
      .d(input_layer[152]),
      .e(~input_layer[1151]),
      .y(Y[900]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron901_1
  function_5 neuron901_1 (
      .a(input_layer[1303]),
      .b(input_layer[115]),
      .y(Y[901]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron902_1
  function_117 neuron902_1 (
      .a(~input_layer[1945]),
      .b(~input_layer[984]),
      .c(input_layer[108]),
      .d(~input_layer[1964]),
      .e(input_layer[391]),
      .f(~input_layer[2028]),
      .y(Y[902]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron903_1
  function_167 neuron903_1 (
      .a(input_layer[1467]),
      .b(~input_layer[1709]),
      .c(input_layer[2217]),
      .d(~input_layer[1826]),
      .e(~input_layer[674]),
      .y(Y[903]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron904_1
  function_40 neuron904_1 (
      .a(~input_layer[1624]),
      .b(input_layer[1308]),
      .c(~input_layer[542]),
      .d(~input_layer[629]),
      .e(~input_layer[1745]),
      .f(~input_layer[998]),
      .y(Y[904]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron905_1
  function_48 neuron905_1 (
      .a(input_layer[279]),
      .b(~input_layer[820]),
      .c(input_layer[142]),
      .d(~input_layer[699]),
      .e(~input_layer[1814]),
      .y(Y[905]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron906_1
  function_30 neuron906_1 (
      .a(input_layer[513]),
      .b(~input_layer[1917]),
      .c(~input_layer[1569]),
      .d(~input_layer[1644]),
      .y(Y[906]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron907_1
  function_248 neuron907_1 (
      .a(~input_layer[552]),
      .b(input_layer[205]),
      .c(~input_layer[1956]),
      .d(~input_layer[2215]),
      .e(input_layer[1539]),
      .f(~input_layer[1260]),
      .y(Y[907]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron908_1
  function_21 neuron908_1 (
      .a(~input_layer[1157]),
      .b(~input_layer[1073]),
      .c(input_layer[1618]),
      .d(input_layer[450]),
      .y(Y[908]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron909_1
  function_183 neuron909_1 (
      .a(input_layer[803]),
      .b(~input_layer[894]),
      .c(input_layer[1907]),
      .d(input_layer[1567]),
      .e(input_layer[416]),
      .f(~input_layer[1975]),
      .y(Y[909]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron910_1
  function_18 neuron910_1 (
      .a(~input_layer[359]),
      .b(~input_layer[2002]),
      .c(~input_layer[1340]),
      .d(~input_layer[1198]),
      .e(~input_layer[2088]),
      .y(Y[910]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_284 for neuron911_1
  function_284 neuron911_1 (
      .a(~input_layer[1549]),
      .b(input_layer[1964]),
      .c(~input_layer[926]),
      .d(input_layer[398]),
      .e(input_layer[1407]),
      .f(~input_layer[1382]),
      .y(Y[911]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron912_1
  function_125 neuron912_1 (
      .a(~input_layer[2164]),
      .b(input_layer[1826]),
      .c(~input_layer[2056]),
      .d(~input_layer[1767]),
      .e(~input_layer[2328]),
      .y(Y[912]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron913_1
  function_54 neuron913_1 (
      .a(input_layer[1729]),
      .b(input_layer[1195]),
      .c(input_layer[199]),
      .d(input_layer[788]),
      .e(input_layer[1951]),
      .f(input_layer[1601]),
      .y(Y[913]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron914_1
  function_35 neuron914_1 (
      .a(~input_layer[1024]),
      .b(input_layer[1047]),
      .c(~input_layer[861]),
      .d(~input_layer[684]),
      .e(input_layer[37]),
      .y(Y[914]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron915_1
  function_60 neuron915_1 (
      .a(~input_layer[317]),
      .b(input_layer[811]),
      .c(~input_layer[184]),
      .d(~input_layer[204]),
      .e(~input_layer[1264]),
      .f(~input_layer[593]),
      .y(Y[915]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron916_1
  function_107 neuron916_1 (
      .a(~input_layer[478]),
      .b(input_layer[1318]),
      .c(~input_layer[352]),
      .d(~input_layer[673]),
      .y(Y[916]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron917_1
  function_3 neuron917_1 (
      .a(input_layer[1211]),
      .b(input_layer[488]),
      .c(input_layer[358]),
      .d(~input_layer[1193]),
      .e(input_layer[1403]),
      .y(Y[917]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_285 for neuron918_1
  function_285 neuron918_1 (
      .a(~input_layer[1142]),
      .b(input_layer[2057]),
      .c(input_layer[1425]),
      .d(~input_layer[1459]),
      .e(~input_layer[1557]),
      .f(~input_layer[2258]),
      .y(Y[918]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron919_1
  function_107 neuron919_1 (
      .a(~input_layer[296]),
      .b(~input_layer[670]),
      .c(input_layer[886]),
      .d(input_layer[930]),
      .y(Y[919]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron920_1
  function_28 neuron920_1 (
      .a(input_layer[742]),
      .b(input_layer[2000]),
      .c(~input_layer[1053]),
      .d(input_layer[1234]),
      .e(input_layer[1782]),
      .f(~input_layer[120]),
      .y(Y[920]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron921_1
  function_128 neuron921_1 (
      .a(~input_layer[1893]),
      .b(input_layer[361]),
      .c(~input_layer[1910]),
      .d(~input_layer[340]),
      .y(Y[921]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_280 for neuron922_1
  function_280 neuron922_1 (
      .a(input_layer[2124]),
      .b(input_layer[431]),
      .c(input_layer[577]),
      .d(~input_layer[819]),
      .e(input_layer[732]),
      .f(input_layer[1573]),
      .y(Y[922]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron923_1
  function_286 neuron923_1 (
      .a(~input_layer[1212]),
      .b(~input_layer[1292]),
      .c(input_layer[2282]),
      .d(input_layer[110]),
      .e(input_layer[626]),
      .y(Y[923]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_250 for neuron924_1
  function_250 neuron924_1 (
      .a(input_layer[746]),
      .b(~input_layer[1564]),
      .c(input_layer[1003]),
      .d(input_layer[1642]),
      .e(input_layer[397]),
      .f(~input_layer[1335]),
      .y(Y[924]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron925_1
  function_34 neuron925_1 (
      .a(input_layer[1327]),
      .b(~input_layer[748]),
      .c(input_layer[2308]),
      .d(input_layer[2022]),
      .e(~input_layer[1034]),
      .y(Y[925]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_287 for neuron926_1
  function_287 neuron926_1 (
      .a(~input_layer[133]),
      .b(~input_layer[1939]),
      .c(input_layer[825]),
      .d(input_layer[709]),
      .e(~input_layer[1536]),
      .f(~input_layer[1813]),
      .y(Y[926]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_288 for neuron927_1
  function_288 neuron927_1 (
      .a(~input_layer[1366]),
      .b(input_layer[1860]),
      .c(~input_layer[1636]),
      .d(input_layer[1938]),
      .e(input_layer[2051]),
      .f(~input_layer[265]),
      .y(Y[927]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron928_1
  function_65 neuron928_1 (
      .a(~input_layer[898]),
      .b(~input_layer[2034]),
      .c(~input_layer[438]),
      .d(input_layer[1375]),
      .e(~input_layer[1511]),
      .f(input_layer[103]),
      .y(Y[928]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron929_1
  function_146 neuron929_1 (
      .a(input_layer[213]),
      .b(input_layer[2335]),
      .c(~input_layer[1893]),
      .d(input_layer[2258]),
      .e(~input_layer[916]),
      .y(Y[929]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_289 for neuron930_1
  function_289 neuron930_1 (
      .a(~input_layer[723]),
      .b(~input_layer[1841]),
      .c(input_layer[498]),
      .d(input_layer[1939]),
      .e(~input_layer[1281]),
      .f(input_layer[2099]),
      .y(Y[930]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron931_1
  function_125 neuron931_1 (
      .a(input_layer[949]),
      .b(~input_layer[1461]),
      .c(~input_layer[1708]),
      .d(~input_layer[272]),
      .e(~input_layer[68]),
      .y(Y[931]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron932_1
  function_52 neuron932_1 (
      .a(~input_layer[467]),
      .b(input_layer[1280]),
      .c(~input_layer[690]),
      .d(input_layer[1878]),
      .e(~input_layer[1450]),
      .y(Y[932]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron933_1
  function_116 neuron933_1 (
      .a(input_layer[1913]),
      .b(~input_layer[1707]),
      .c(input_layer[558]),
      .d(input_layer[1061]),
      .y(Y[933]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron934_1
  function_11 neuron934_1 (
      .a(input_layer[364]),
      .b(input_layer[133]),
      .c(~input_layer[1452]),
      .d(input_layer[131]),
      .y(Y[934]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron935_1
  function_290 neuron935_1 (
      .a(~input_layer[981]),
      .b(input_layer[1405]),
      .c(input_layer[565]),
      .d(~input_layer[1758]),
      .e(~input_layer[470]),
      .y(Y[935]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron936_1
  function_125 neuron936_1 (
      .a(input_layer[654]),
      .b(~input_layer[730]),
      .c(~input_layer[2296]),
      .d(~input_layer[2171]),
      .e(input_layer[461]),
      .y(Y[936]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_262 for neuron937_1
  function_262 neuron937_1 (
      .a(input_layer[1156]),
      .b(input_layer[2241]),
      .c(input_layer[1427]),
      .d(input_layer[2270]),
      .e(input_layer[0]),
      .f(input_layer[153]),
      .y(Y[937]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_291 for neuron938_1
  function_291 neuron938_1 (
      .a(~input_layer[1495]),
      .b(~input_layer[1784]),
      .c(input_layer[2202]),
      .d(~input_layer[1259]),
      .e(input_layer[145]),
      .f(input_layer[480]),
      .y(Y[938]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron939_1
  function_12 neuron939_1 (
      .a(~input_layer[1504]),
      .b(input_layer[1314]),
      .c(~input_layer[1712]),
      .y(Y[939]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron940_1
  function_49 neuron940_1 (
      .a(input_layer[822]),
      .b(input_layer[2239]),
      .c(input_layer[394]),
      .d(input_layer[405]),
      .e(~input_layer[287]),
      .f(~input_layer[1533]),
      .y(Y[940]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_292 for neuron941_1
  function_292 neuron941_1 (
      .a(input_layer[1496]),
      .b(~input_layer[2115]),
      .c(~input_layer[682]),
      .d(~input_layer[138]),
      .e(~input_layer[2286]),
      .f(input_layer[1781]),
      .y(Y[941]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron942_1
  function_26 neuron942_1 (
      .a(~input_layer[192]),
      .b(~input_layer[375]),
      .y(Y[942]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron943_1
  function_44 neuron943_1 (
      .a(~input_layer[364]),
      .b(input_layer[808]),
      .c(input_layer[643]),
      .y(Y[943]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron944_1
  function_5 neuron944_1 (
      .a(input_layer[1417]),
      .b(~input_layer[1866]),
      .y(Y[944]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_293 for neuron945_1
  function_293 neuron945_1 (
      .a(input_layer[1453]),
      .b(input_layer[1365]),
      .c(~input_layer[1412]),
      .d(input_layer[986]),
      .e(~input_layer[1678]),
      .f(input_layer[622]),
      .y(Y[945]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron946_1
  function_100 neuron946_1 (
      .a(input_layer[1373]),
      .b(input_layer[1065]),
      .c(~input_layer[899]),
      .y(Y[946]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron947_1
  function_45 neuron947_1 (
      .a(~input_layer[310]),
      .b(~input_layer[432]),
      .c(~input_layer[1675]),
      .d(input_layer[625]),
      .e(~input_layer[2232]),
      .f(input_layer[485]),
      .y(Y[947]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_160 for neuron948_1
  function_160 neuron948_1 (
      .a(input_layer[231]),
      .b(~input_layer[1612]),
      .c(~input_layer[1710]),
      .d(~input_layer[535]),
      .e(~input_layer[376]),
      .y(Y[948]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron949_1
  function_286 neuron949_1 (
      .a(~input_layer[1620]),
      .b(input_layer[617]),
      .c(~input_layer[621]),
      .d(~input_layer[472]),
      .e(input_layer[2177]),
      .y(Y[949]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron950_1
  function_12 neuron950_1 (
      .a(~input_layer[2137]),
      .b(~input_layer[1315]),
      .c(~input_layer[1666]),
      .y(Y[950]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_294 for neuron951_1
  function_294 neuron951_1 (
      .a(input_layer[886]),
      .b(~input_layer[2204]),
      .c(~input_layer[1368]),
      .d(input_layer[1985]),
      .e(~input_layer[2336]),
      .f(~input_layer[981]),
      .y(Y[951]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron952_1
  function_16 neuron952_1 (
      .a(input_layer[2318]),
      .b(input_layer[2115]),
      .c(input_layer[1141]),
      .y(Y[952]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron953_1
  function_91 neuron953_1 (
      .a(input_layer[1778]),
      .b(input_layer[2326]),
      .c(input_layer[1313]),
      .d(~input_layer[240]),
      .e(~input_layer[2183]),
      .f(input_layer[2104]),
      .y(Y[953]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_295 for neuron954_1
  function_295 neuron954_1 (
      .a(~input_layer[1278]),
      .b(input_layer[1266]),
      .c(input_layer[1211]),
      .d(input_layer[757]),
      .e(input_layer[1804]),
      .f(~input_layer[253]),
      .y(Y[954]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_296 for neuron955_1
  function_296 neuron955_1 (
      .a(~input_layer[198]),
      .b(~input_layer[2236]),
      .c(~input_layer[1033]),
      .d(input_layer[1602]),
      .e(input_layer[1940]),
      .f(~input_layer[907]),
      .y(Y[955]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron956_1
  function_10 neuron956_1 (
      .a(input_layer[1988]),
      .b(~input_layer[974]),
      .c(~input_layer[729]),
      .d(input_layer[979]),
      .y(Y[956]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron957_1
  function_11 neuron957_1 (
      .a(input_layer[1190]),
      .b(input_layer[406]),
      .c(input_layer[1842]),
      .d(~input_layer[967]),
      .y(Y[957]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron958_1
  function_24 neuron958_1 (
      .a(input_layer[491]),
      .y(Y[958]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron959_1
  function_210 neuron959_1 (
      .a(~input_layer[1131]),
      .b(input_layer[287]),
      .c(input_layer[1943]),
      .d(~input_layer[552]),
      .e(input_layer[1821]),
      .y(Y[959]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron960_1
  function_95 neuron960_1 (
      .a(input_layer[2077]),
      .b(~input_layer[1453]),
      .c(input_layer[553]),
      .d(~input_layer[608]),
      .y(Y[960]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_297 for neuron961_1
  function_297 neuron961_1 (
      .a(~input_layer[839]),
      .b(input_layer[1035]),
      .c(input_layer[947]),
      .d(~input_layer[2212]),
      .e(~input_layer[2047]),
      .y(Y[961]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron962_1
  function_162 neuron962_1 (
      .a(~input_layer[2073]),
      .b(~input_layer[227]),
      .c(input_layer[966]),
      .d(input_layer[1480]),
      .e(input_layer[2107]),
      .y(Y[962]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron963_1
  function_298 neuron963_1 (
      .a(~input_layer[1654]),
      .b(input_layer[1604]),
      .c(input_layer[517]),
      .d(~input_layer[1816]),
      .e(~input_layer[1023]),
      .y(Y[963]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron964_1
  function_16 neuron964_1 (
      .a(input_layer[2326]),
      .b(~input_layer[555]),
      .c(~input_layer[1056]),
      .y(Y[964]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron965_1
  function_299 neuron965_1 (
      .a(input_layer[1383]),
      .b(input_layer[1335]),
      .c(~input_layer[912]),
      .d(input_layer[404]),
      .e(input_layer[1364]),
      .f(input_layer[1476]),
      .y(Y[965]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron966_1
  function_76 neuron966_1 (
      .a(~input_layer[1243]),
      .b(~input_layer[2209]),
      .c(~input_layer[2310]),
      .d(~input_layer[1769]),
      .e(~input_layer[2292]),
      .f(~input_layer[1852]),
      .y(Y[966]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_300 for neuron967_1
  function_300 neuron967_1 (
      .a(input_layer[1629]),
      .b(input_layer[1255]),
      .c(input_layer[1863]),
      .d(~input_layer[937]),
      .e(~input_layer[1822]),
      .y(Y[967]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron968_1
  function_149 neuron968_1 (
      .a(~input_layer[394]),
      .b(~input_layer[1149]),
      .c(~input_layer[1490]),
      .d(input_layer[1907]),
      .y(Y[968]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron969_1
  function_210 neuron969_1 (
      .a(input_layer[958]),
      .b(~input_layer[373]),
      .c(input_layer[2324]),
      .d(input_layer[1424]),
      .e(input_layer[488]),
      .y(Y[969]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron970_1
  function_64 neuron970_1 (
      .a(input_layer[1785]),
      .b(input_layer[451]),
      .c(~input_layer[1802]),
      .d(input_layer[1089]),
      .e(input_layer[713]),
      .y(Y[970]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron971_1
  function_146 neuron971_1 (
      .a(input_layer[916]),
      .b(input_layer[1856]),
      .c(input_layer[633]),
      .d(~input_layer[1710]),
      .e(input_layer[733]),
      .y(Y[971]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_301 for neuron972_1
  function_301 neuron972_1 (
      .a(~input_layer[2133]),
      .b(input_layer[1840]),
      .c(~input_layer[669]),
      .d(~input_layer[1482]),
      .e(input_layer[1783]),
      .f(input_layer[937]),
      .y(Y[972]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_302 for neuron973_1
  function_302 neuron973_1 (
      .a(~input_layer[575]),
      .b(input_layer[1168]),
      .c(input_layer[1842]),
      .d(input_layer[1880]),
      .e(~input_layer[1995]),
      .y(Y[973]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron974_1
  function_107 neuron974_1 (
      .a(~input_layer[1634]),
      .b(~input_layer[1627]),
      .c(~input_layer[1836]),
      .d(~input_layer[1200]),
      .y(Y[974]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron975_1
  function_25 neuron975_1 (
      .a(input_layer[1107]),
      .b(input_layer[2080]),
      .c(input_layer[1170]),
      .d(~input_layer[1629]),
      .e(input_layer[431]),
      .y(Y[975]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron976_1
  function_11 neuron976_1 (
      .a(input_layer[663]),
      .b(input_layer[752]),
      .c(input_layer[1358]),
      .d(input_layer[1371]),
      .y(Y[976]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_174 for neuron977_1
  function_174 neuron977_1 (
      .a(~input_layer[1712]),
      .b(~input_layer[1506]),
      .c(input_layer[806]),
      .d(~input_layer[384]),
      .e(~input_layer[1787]),
      .f(input_layer[773]),
      .y(Y[977]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron978_1
  function_303 neuron978_1 (
      .a(input_layer[1016]),
      .b(input_layer[1796]),
      .c(input_layer[1494]),
      .d(input_layer[822]),
      .e(~input_layer[2221]),
      .f(input_layer[191]),
      .y(Y[978]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron979_1
  function_0 neuron979_1 (
      .a(input_layer[316]),
      .b(~input_layer[546]),
      .c(input_layer[1724]),
      .d(input_layer[1730]),
      .e(input_layer[1819]),
      .y(Y[979]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron980_1
  function_56 neuron980_1 (
      .a(~input_layer[650]),
      .b(input_layer[1546]),
      .c(~input_layer[1908]),
      .d(~input_layer[902]),
      .e(input_layer[1032]),
      .y(Y[980]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron981_1
  function_12 neuron981_1 (
      .a(~input_layer[1944]),
      .b(~input_layer[1737]),
      .c(~input_layer[1776]),
      .y(Y[981]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron982_1
  function_148 neuron982_1 (
      .a(~input_layer[1380]),
      .b(input_layer[1885]),
      .c(~input_layer[146]),
      .d(~input_layer[2332]),
      .y(Y[982]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron983_1
  function_63 neuron983_1 (
      .a(input_layer[2239]),
      .b(input_layer[646]),
      .c(~input_layer[2115]),
      .d(input_layer[818]),
      .y(Y[983]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron984_1
  function_3 neuron984_1 (
      .a(input_layer[1054]),
      .b(input_layer[356]),
      .c(input_layer[1003]),
      .d(~input_layer[792]),
      .e(~input_layer[2199]),
      .y(Y[984]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron985_1
  function_12 neuron985_1 (
      .a(~input_layer[1320]),
      .b(~input_layer[2220]),
      .c(~input_layer[930]),
      .y(Y[985]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron986_1
  function_139 neuron986_1 (
      .a(~input_layer[708]),
      .b(~input_layer[1918]),
      .c(input_layer[569]),
      .d(input_layer[2259]),
      .e(input_layer[2284]),
      .y(Y[986]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron987_1
  function_87 neuron987_1 (
      .a(input_layer[2134]),
      .b(input_layer[2208]),
      .c(input_layer[1520]),
      .d(~input_layer[116]),
      .e(input_layer[2090]),
      .f(input_layer[597]),
      .y(Y[987]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron988_1
  function_248 neuron988_1 (
      .a(~input_layer[1462]),
      .b(~input_layer[790]),
      .c(~input_layer[191]),
      .d(input_layer[475]),
      .e(input_layer[640]),
      .f(input_layer[258]),
      .y(Y[988]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron989_1
  function_43 neuron989_1 (
      .a(input_layer[747]),
      .b(~input_layer[801]),
      .c(~input_layer[1256]),
      .d(~input_layer[2254]),
      .e(~input_layer[1099]),
      .y(Y[989]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_225 for neuron990_1
  function_225 neuron990_1 (
      .a(~input_layer[1460]),
      .b(~input_layer[2326]),
      .c(input_layer[1818]),
      .d(input_layer[969]),
      .e(input_layer[1594]),
      .f(~input_layer[80]),
      .y(Y[990]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_304 for neuron991_1
  function_304 neuron991_1 (
      .a(input_layer[610]),
      .b(~input_layer[1246]),
      .c(~input_layer[322]),
      .d(input_layer[999]),
      .e(~input_layer[2304]),
      .f(input_layer[84]),
      .y(Y[991]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron992_1
  function_181 neuron992_1 (
      .a(~input_layer[2296]),
      .b(input_layer[1198]),
      .c(~input_layer[744]),
      .d(~input_layer[2233]),
      .e(~input_layer[2022]),
      .f(~input_layer[2096]),
      .y(Y[992]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron993_1
  function_99 neuron993_1 (
      .a(input_layer[980]),
      .b(input_layer[2235]),
      .c(~input_layer[1059]),
      .d(input_layer[446]),
      .e(input_layer[393]),
      .f(~input_layer[2263]),
      .y(Y[993]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron994_1
  function_3 neuron994_1 (
      .a(input_layer[1496]),
      .b(input_layer[2224]),
      .c(input_layer[639]),
      .d(input_layer[190]),
      .e(~input_layer[694]),
      .y(Y[994]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron995_1
  function_0 neuron995_1 (
      .a(input_layer[1213]),
      .b(input_layer[1833]),
      .c(~input_layer[724]),
      .d(input_layer[830]),
      .e(~input_layer[1411]),
      .y(Y[995]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron996_1
  function_10 neuron996_1 (
      .a(input_layer[655]),
      .b(~input_layer[2226]),
      .c(input_layer[2115]),
      .d(input_layer[242]),
      .y(Y[996]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron997_1
  function_21 neuron997_1 (
      .a(~input_layer[1999]),
      .b(~input_layer[2148]),
      .c(~input_layer[1899]),
      .d(~input_layer[943]),
      .y(Y[997]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_183 for neuron998_1
  function_183 neuron998_1 (
      .a(input_layer[1544]),
      .b(~input_layer[909]),
      .c(input_layer[1426]),
      .d(~input_layer[1511]),
      .e(input_layer[2340]),
      .f(~input_layer[1979]),
      .y(Y[998]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron999_1
  function_16 neuron999_1 (
      .a(input_layer[2075]),
      .b(~input_layer[1583]),
      .c(~input_layer[1459]),
      .y(Y[999]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1000_1
  function_169 neuron1000_1 (
      .a(input_layer[1197]),
      .b(input_layer[2222]),
      .c(input_layer[975]),
      .d(~input_layer[1306]),
      .e(~input_layer[1633]),
      .f(~input_layer[1723]),
      .y(Y[1000]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_305 for neuron1001_1
  function_305 neuron1001_1 (
      .a(input_layer[1724]),
      .b(input_layer[1423]),
      .c(~input_layer[1052]),
      .d(input_layer[2208]),
      .e(~input_layer[1170]),
      .f(input_layer[652]),
      .y(Y[1001]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron1002_1
  function_69 neuron1002_1 (
      .a(input_layer[1075]),
      .b(input_layer[1946]),
      .c(~input_layer[1977]),
      .d(input_layer[1883]),
      .e(~input_layer[1700]),
      .y(Y[1002]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1003_1
  function_100 neuron1003_1 (
      .a(~input_layer[985]),
      .b(~input_layer[448]),
      .c(input_layer[1426]),
      .y(Y[1003]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1004_1
  function_26 neuron1004_1 (
      .a(~input_layer[1225]),
      .b(~input_layer[1278]),
      .y(Y[1004]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_306 for neuron1005_1
  function_306 neuron1005_1 (
      .a(input_layer[1423]),
      .b(input_layer[939]),
      .c(~input_layer[974]),
      .d(input_layer[650]),
      .e(~input_layer[1978]),
      .f(input_layer[1796]),
      .y(Y[1005]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1006_1
  function_63 neuron1006_1 (
      .a(input_layer[1038]),
      .b(input_layer[364]),
      .c(~input_layer[488]),
      .d(~input_layer[109]),
      .y(Y[1006]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_17 for neuron1007_1
  function_17 neuron1007_1 (
      .a(~input_layer[2067]),
      .b(input_layer[1733]),
      .c(~input_layer[327]),
      .d(input_layer[571]),
      .e(~input_layer[2195]),
      .f(~input_layer[1682]),
      .y(Y[1007]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1008_1
  function_49 neuron1008_1 (
      .a(input_layer[1078]),
      .b(input_layer[2129]),
      .c(input_layer[1319]),
      .d(input_layer[1436]),
      .e(input_layer[1775]),
      .f(input_layer[2336]),
      .y(Y[1008]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1009_1
  function_307 neuron1009_1 (
      .a(~input_layer[222]),
      .b(input_layer[1447]),
      .c(~input_layer[804]),
      .d(~input_layer[243]),
      .e(input_layer[1807]),
      .y(Y[1009]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1010_1
  function_3 neuron1010_1 (
      .a(input_layer[526]),
      .b(input_layer[2318]),
      .c(input_layer[2331]),
      .d(~input_layer[1407]),
      .e(input_layer[1822]),
      .y(Y[1010]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1011_1
  function_21 neuron1011_1 (
      .a(~input_layer[1673]),
      .b(~input_layer[1353]),
      .c(~input_layer[1683]),
      .d(~input_layer[1583]),
      .y(Y[1011]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1012] = 1'b0;

  // instantiate function_239 for neuron1013_1
  function_239 neuron1013_1 (
      .a(input_layer[2237]),
      .b(input_layer[948]),
      .c(input_layer[1082]),
      .d(~input_layer[1335]),
      .e(~input_layer[1489]),
      .y(Y[1013]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1014_1
  function_64 neuron1014_1 (
      .a(input_layer[1041]),
      .b(input_layer[2225]),
      .c(input_layer[1289]),
      .d(input_layer[1656]),
      .e(~input_layer[1063]),
      .y(Y[1014]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1015_1
  function_12 neuron1015_1 (
      .a(~input_layer[578]),
      .b(~input_layer[433]),
      .c(~input_layer[734]),
      .y(Y[1015]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1016_1
  function_162 neuron1016_1 (
      .a(~input_layer[2041]),
      .b(~input_layer[309]),
      .c(~input_layer[441]),
      .d(~input_layer[1239]),
      .e(~input_layer[380]),
      .y(Y[1016]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1017_1
  function_4 neuron1017_1 (
      .a(input_layer[2307]),
      .b(~input_layer[1065]),
      .c(~input_layer[1561]),
      .d(input_layer[1064]),
      .e(input_layer[756]),
      .y(Y[1017]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1018_1
  function_21 neuron1018_1 (
      .a(~input_layer[290]),
      .b(input_layer[1286]),
      .c(~input_layer[2086]),
      .d(~input_layer[2331]),
      .y(Y[1018]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1019_1
  function_14 neuron1019_1 (
      .a(~input_layer[543]),
      .b(~input_layer[860]),
      .c(~input_layer[1582]),
      .d(~input_layer[434]),
      .e(~input_layer[1343]),
      .y(Y[1019]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1020_1
  function_21 neuron1020_1 (
      .a(~input_layer[616]),
      .b(~input_layer[1437]),
      .c(input_layer[970]),
      .d(~input_layer[538]),
      .y(Y[1020]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1021_1
  function_3 neuron1021_1 (
      .a(input_layer[995]),
      .b(input_layer[2237]),
      .c(input_layer[222]),
      .d(~input_layer[651]),
      .e(input_layer[1605]),
      .y(Y[1021]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1022_1
  function_63 neuron1022_1 (
      .a(input_layer[949]),
      .b(input_layer[871]),
      .c(~input_layer[681]),
      .d(~input_layer[1635]),
      .y(Y[1022]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1023_1
  function_92 neuron1023_1 (
      .a(input_layer[798]),
      .b(input_layer[2127]),
      .c(input_layer[348]),
      .d(~input_layer[1211]),
      .y(Y[1023]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1024_1
  function_1 neuron1024_1 (
      .a(~input_layer[1660]),
      .b(~input_layer[357]),
      .c(~input_layer[1781]),
      .d(~input_layer[1290]),
      .e(input_layer[524]),
      .f(input_layer[1400]),
      .y(Y[1024]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1025_1
  function_32 neuron1025_1 (
      .a(input_layer[1069]),
      .b(input_layer[1360]),
      .c(~input_layer[1478]),
      .d(~input_layer[585]),
      .y(Y[1025]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_280 for neuron1026_1
  function_280 neuron1026_1 (
      .a(input_layer[1999]),
      .b(input_layer[366]),
      .c(input_layer[120]),
      .d(~input_layer[2318]),
      .e(~input_layer[1487]),
      .f(input_layer[243]),
      .y(Y[1026]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1027_1
  function_167 neuron1027_1 (
      .a(~input_layer[2141]),
      .b(input_layer[641]),
      .c(~input_layer[1488]),
      .d(~input_layer[1893]),
      .e(input_layer[1298]),
      .y(Y[1027]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1028_1
  function_181 neuron1028_1 (
      .a(~input_layer[203]),
      .b(~input_layer[809]),
      .c(~input_layer[439]),
      .d(~input_layer[1559]),
      .e(~input_layer[2140]),
      .f(input_layer[879]),
      .y(Y[1028]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1029_1
  function_44 neuron1029_1 (
      .a(input_layer[1300]),
      .b(~input_layer[1245]),
      .c(~input_layer[1718]),
      .y(Y[1029]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_308 for neuron1030_1
  function_308 neuron1030_1 (
      .a(input_layer[654]),
      .b(~input_layer[1911]),
      .c(input_layer[1331]),
      .d(input_layer[818]),
      .e(~input_layer[1808]),
      .f(~input_layer[118]),
      .y(Y[1030]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1031_1
  function_53 neuron1031_1 (
      .a(input_layer[212]),
      .b(input_layer[1579]),
      .c(~input_layer[2299]),
      .d(input_layer[869]),
      .e(input_layer[722]),
      .y(Y[1031]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1032_1
  function_25 neuron1032_1 (
      .a(input_layer[836]),
      .b(input_layer[587]),
      .c(~input_layer[970]),
      .d(input_layer[1341]),
      .e(~input_layer[888]),
      .y(Y[1032]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1033_1
  function_56 neuron1033_1 (
      .a(~input_layer[2142]),
      .b(~input_layer[2002]),
      .c(input_layer[405]),
      .d(input_layer[1294]),
      .e(~input_layer[1873]),
      .y(Y[1033]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1034_1
  function_14 neuron1034_1 (
      .a(~input_layer[1389]),
      .b(~input_layer[1422]),
      .c(~input_layer[585]),
      .d(~input_layer[449]),
      .e(~input_layer[564]),
      .y(Y[1034]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1035_1
  function_162 neuron1035_1 (
      .a(~input_layer[1605]),
      .b(~input_layer[552]),
      .c(~input_layer[2249]),
      .d(~input_layer[1315]),
      .e(input_layer[1654]),
      .y(Y[1035]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1036_1
  function_12 neuron1036_1 (
      .a(~input_layer[581]),
      .b(~input_layer[836]),
      .c(~input_layer[1899]),
      .y(Y[1036]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1037_1
  function_31 neuron1037_1 (
      .a(input_layer[1586]),
      .b(input_layer[440]),
      .c(input_layer[230]),
      .d(input_layer[1167]),
      .e(input_layer[515]),
      .f(input_layer[755]),
      .y(Y[1037]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_309 for neuron1038_1
  function_309 neuron1038_1 (
      .a(input_layer[760]),
      .b(~input_layer[863]),
      .c(~input_layer[1417]),
      .d(input_layer[623]),
      .e(~input_layer[561]),
      .f(~input_layer[984]),
      .y(Y[1038]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1039_1
  function_25 neuron1039_1 (
      .a(input_layer[296]),
      .b(input_layer[1505]),
      .c(input_layer[2218]),
      .d(input_layer[718]),
      .e(input_layer[2305]),
      .y(Y[1039]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_136 for neuron1040_1
  function_136 neuron1040_1 (
      .a(input_layer[203]),
      .b(~input_layer[1754]),
      .c(~input_layer[1648]),
      .d(input_layer[696]),
      .e(~input_layer[295]),
      .f(input_layer[2259]),
      .y(Y[1040]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_291 for neuron1041_1
  function_291 neuron1041_1 (
      .a(~input_layer[1305]),
      .b(input_layer[1015]),
      .c(~input_layer[1918]),
      .d(~input_layer[2313]),
      .e(~input_layer[310]),
      .f(input_layer[925]),
      .y(Y[1041]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1042_1
  function_4 neuron1042_1 (
      .a(input_layer[1246]),
      .b(input_layer[238]),
      .c(input_layer[315]),
      .d(~input_layer[1104]),
      .e(~input_layer[788]),
      .y(Y[1042]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1043_1
  function_67 neuron1043_1 (
      .a(input_layer[1198]),
      .b(input_layer[430]),
      .c(~input_layer[1639]),
      .d(input_layer[1565]),
      .e(input_layer[339]),
      .y(Y[1043]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1044_1
  function_12 neuron1044_1 (
      .a(~input_layer[1145]),
      .b(~input_layer[2002]),
      .c(input_layer[1195]),
      .y(Y[1044]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1045_1
  function_76 neuron1045_1 (
      .a(~input_layer[1887]),
      .b(~input_layer[1417]),
      .c(~input_layer[498]),
      .d(~input_layer[244]),
      .e(~input_layer[755]),
      .f(~input_layer[2091]),
      .y(Y[1045]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1046_1
  function_14 neuron1046_1 (
      .a(~input_layer[835]),
      .b(~input_layer[1168]),
      .c(input_layer[573]),
      .d(~input_layer[1669]),
      .e(input_layer[606]),
      .y(Y[1046]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1047_1
  function_125 neuron1047_1 (
      .a(~input_layer[1087]),
      .b(~input_layer[1321]),
      .c(~input_layer[2077]),
      .d(input_layer[1356]),
      .e(~input_layer[1849]),
      .y(Y[1047]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1048_1
  function_5 neuron1048_1 (
      .a(input_layer[875]),
      .b(input_layer[2226]),
      .y(Y[1048]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_310 for neuron1049_1
  function_310 neuron1049_1 (
      .a(~input_layer[1419]),
      .b(input_layer[1313]),
      .c(input_layer[1235]),
      .d(~input_layer[816]),
      .e(input_layer[324]),
      .f(~input_layer[676]),
      .y(Y[1049]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron1050_1
  function_115 neuron1050_1 (
      .a(input_layer[1544]),
      .b(~input_layer[307]),
      .c(input_layer[785]),
      .d(input_layer[1254]),
      .e(~input_layer[1732]),
      .y(Y[1050]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_311 for neuron1051_1
  function_311 neuron1051_1 (
      .a(~input_layer[1169]),
      .b(input_layer[1942]),
      .c(input_layer[1787]),
      .d(input_layer[703]),
      .e(input_layer[1854]),
      .f(input_layer[1320]),
      .y(Y[1051]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron1052_1
  function_130 neuron1052_1 (
      .a(input_layer[819]),
      .b(input_layer[285]),
      .c(input_layer[979]),
      .d(~input_layer[2253]),
      .e(~input_layer[1163]),
      .f(input_layer[710]),
      .y(Y[1052]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_312 for neuron1053_1
  function_312 neuron1053_1 (
      .a(input_layer[1051]),
      .b(input_layer[317]),
      .c(~input_layer[1510]),
      .d(~input_layer[470]),
      .e(~input_layer[896]),
      .f(input_layer[1850]),
      .y(Y[1053]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1054_1
  function_67 neuron1054_1 (
      .a(input_layer[1578]),
      .b(~input_layer[2159]),
      .c(input_layer[1837]),
      .d(input_layer[2309]),
      .e(input_layer[1302]),
      .y(Y[1054]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1055_1
  function_95 neuron1055_1 (
      .a(~input_layer[1888]),
      .b(input_layer[2211]),
      .c(~input_layer[2153]),
      .d(input_layer[2084]),
      .y(Y[1055]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1056_1
  function_16 neuron1056_1 (
      .a(input_layer[783]),
      .b(input_layer[745]),
      .c(~input_layer[1491]),
      .y(Y[1056]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_313 for neuron1057_1
  function_313 neuron1057_1 (
      .a(input_layer[1044]),
      .b(~input_layer[2288]),
      .c(~input_layer[2032]),
      .d(input_layer[322]),
      .e(~input_layer[1345]),
      .f(~input_layer[1620]),
      .y(Y[1057]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1058_1
  function_188 neuron1058_1 (
      .a(input_layer[1300]),
      .b(input_layer[1339]),
      .c(~input_layer[410]),
      .d(input_layer[1666]),
      .e(~input_layer[1239]),
      .f(input_layer[240]),
      .y(Y[1058]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1059_1
  function_16 neuron1059_1 (
      .a(input_layer[1000]),
      .b(input_layer[275]),
      .c(~input_layer[1392]),
      .y(Y[1059]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_314 for neuron1060_1
  function_314 neuron1060_1 (
      .a(input_layer[912]),
      .b(~input_layer[284]),
      .c(~input_layer[979]),
      .d(~input_layer[289]),
      .e(~input_layer[1378]),
      .f(input_layer[248]),
      .y(Y[1060]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1061_1
  function_32 neuron1061_1 (
      .a(~input_layer[377]),
      .b(input_layer[763]),
      .c(input_layer[1328]),
      .d(input_layer[416]),
      .y(Y[1061]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1062_1
  function_4 neuron1062_1 (
      .a(input_layer[454]),
      .b(~input_layer[268]),
      .c(input_layer[2022]),
      .d(input_layer[1790]),
      .e(input_layer[1823]),
      .y(Y[1062]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_30 for neuron1063_1
  function_30 neuron1063_1 (
      .a(input_layer[311]),
      .b(input_layer[118]),
      .c(~input_layer[1648]),
      .d(~input_layer[687]),
      .y(Y[1063]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_82 for neuron1064_1
  function_82 neuron1064_1 (
      .a(~input_layer[2234]),
      .b(~input_layer[2204]),
      .c(input_layer[1168]),
      .d(input_layer[1675]),
      .e(~input_layer[1989]),
      .y(Y[1064]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1065_1
  function_307 neuron1065_1 (
      .a(~input_layer[714]),
      .b(~input_layer[314]),
      .c(input_layer[1548]),
      .d(~input_layer[1830]),
      .e(~input_layer[710]),
      .y(Y[1065]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_315 for neuron1066_1
  function_315 neuron1066_1 (
      .a(input_layer[2090]),
      .b(~input_layer[2316]),
      .c(~input_layer[893]),
      .d(input_layer[415]),
      .e(~input_layer[1268]),
      .f(~input_layer[1009]),
      .y(Y[1066]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1067_1
  function_162 neuron1067_1 (
      .a(~input_layer[494]),
      .b(~input_layer[431]),
      .c(input_layer[950]),
      .d(~input_layer[2110]),
      .e(~input_layer[1584]),
      .y(Y[1067]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_109 for neuron1068_1
  function_109 neuron1068_1 (
      .a(input_layer[2216]),
      .b(~input_layer[1212]),
      .c(input_layer[818]),
      .d(input_layer[1072]),
      .e(~input_layer[665]),
      .f(input_layer[1067]),
      .y(Y[1068]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1069_1
  function_44 neuron1069_1 (
      .a(~input_layer[548]),
      .b(input_layer[1107]),
      .c(~input_layer[829]),
      .y(Y[1069]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1070_1
  function_12 neuron1070_1 (
      .a(~input_layer[1583]),
      .b(~input_layer[1360]),
      .c(input_layer[854]),
      .y(Y[1070]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1071_1
  function_12 neuron1071_1 (
      .a(~input_layer[565]),
      .b(~input_layer[1670]),
      .c(input_layer[618]),
      .y(Y[1071]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_316 for neuron1072_1
  function_316 neuron1072_1 (
      .a(input_layer[595]),
      .b(~input_layer[1971]),
      .c(input_layer[1758]),
      .d(input_layer[1994]),
      .e(input_layer[2334]),
      .f(input_layer[1867]),
      .y(Y[1072]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1073_1
  function_12 neuron1073_1 (
      .a(~input_layer[2290]),
      .b(~input_layer[694]),
      .c(~input_layer[242]),
      .y(Y[1073]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_317 for neuron1074_1
  function_317 neuron1074_1 (
      .a(~input_layer[1701]),
      .b(input_layer[487]),
      .c(~input_layer[434]),
      .d(~input_layer[1166]),
      .e(~input_layer[1433]),
      .f(~input_layer[1612]),
      .y(Y[1074]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_290 for neuron1075_1
  function_290 neuron1075_1 (
      .a(~input_layer[661]),
      .b(~input_layer[104]),
      .c(input_layer[2237]),
      .d(input_layer[2149]),
      .e(~input_layer[1049]),
      .y(Y[1075]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1076] = 1'b1;

  // instantiate function_307 for neuron1077_1
  function_307 neuron1077_1 (
      .a(~input_layer[450]),
      .b(input_layer[817]),
      .c(input_layer[804]),
      .d(~input_layer[2023]),
      .e(~input_layer[883]),
      .y(Y[1077]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_318 for neuron1078_1
  function_318 neuron1078_1 (
      .a(~input_layer[780]),
      .b(input_layer[1350]),
      .c(~input_layer[1065]),
      .d(input_layer[38]),
      .e(~input_layer[1090]),
      .f(~input_layer[83]),
      .y(Y[1078]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1079_1
  function_24 neuron1079_1 (
      .a(~input_layer[2133]),
      .y(Y[1079]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1080_1
  function_26 neuron1080_1 (
      .a(~input_layer[2220]),
      .b(input_layer[1480]),
      .y(Y[1080]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1081_1
  function_319 neuron1081_1 (
      .a(input_layer[707]),
      .b(input_layer[1967]),
      .c(~input_layer[1394]),
      .d(input_layer[557]),
      .e(input_layer[1887]),
      .f(~input_layer[1198]),
      .y(Y[1081]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1082_1
  function_11 neuron1082_1 (
      .a(input_layer[886]),
      .b(input_layer[598]),
      .c(input_layer[516]),
      .d(~input_layer[1401]),
      .y(Y[1082]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1083_1
  function_107 neuron1083_1 (
      .a(~input_layer[494]),
      .b(input_layer[382]),
      .c(~input_layer[2306]),
      .d(~input_layer[730]),
      .y(Y[1083]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1084_1
  function_44 neuron1084_1 (
      .a(~input_layer[1366]),
      .b(input_layer[966]),
      .c(input_layer[105]),
      .y(Y[1084]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1085_1
  function_21 neuron1085_1 (
      .a(~input_layer[2060]),
      .b(~input_layer[308]),
      .c(~input_layer[219]),
      .d(~input_layer[2043]),
      .y(Y[1085]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_142 for neuron1086_1
  function_142 neuron1086_1 (
      .a(~input_layer[231]),
      .b(input_layer[554]),
      .c(input_layer[717]),
      .d(input_layer[2134]),
      .e(input_layer[630]),
      .y(Y[1086]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1087_1
  function_18 neuron1087_1 (
      .a(~input_layer[1946]),
      .b(~input_layer[2129]),
      .c(input_layer[1488]),
      .d(~input_layer[1687]),
      .e(~input_layer[2319]),
      .y(Y[1087]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1088_1
  function_25 neuron1088_1 (
      .a(input_layer[2073]),
      .b(input_layer[408]),
      .c(input_layer[1602]),
      .d(~input_layer[1575]),
      .e(~input_layer[1561]),
      .y(Y[1088]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1089_1
  function_0 neuron1089_1 (
      .a(input_layer[1741]),
      .b(input_layer[230]),
      .c(input_layer[2083]),
      .d(input_layer[2069]),
      .e(~input_layer[1406]),
      .y(Y[1089]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_194 for neuron1090_1
  function_194 neuron1090_1 (
      .a(input_layer[988]),
      .b(~input_layer[539]),
      .c(input_layer[683]),
      .d(input_layer[428]),
      .e(input_layer[1089]),
      .f(input_layer[2252]),
      .y(Y[1090]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1091_1
  function_12 neuron1091_1 (
      .a(input_layer[1042]),
      .b(~input_layer[1709]),
      .c(~input_layer[2042]),
      .y(Y[1091]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron1092_1
  function_286 neuron1092_1 (
      .a(input_layer[1498]),
      .b(~input_layer[968]),
      .c(input_layer[1793]),
      .d(~input_layer[557]),
      .e(input_layer[47]),
      .y(Y[1092]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_320 for neuron1093_1
  function_320 neuron1093_1 (
      .a(~input_layer[962]),
      .b(input_layer[1838]),
      .c(~input_layer[1134]),
      .d(~input_layer[1270]),
      .e(input_layer[1358]),
      .f(~input_layer[456]),
      .y(Y[1093]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1094_1
  function_104 neuron1094_1 (
      .a(~input_layer[834]),
      .b(input_layer[2207]),
      .c(~input_layer[790]),
      .y(Y[1094]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1095_1
  function_16 neuron1095_1 (
      .a(input_layer[368]),
      .b(~input_layer[883]),
      .c(input_layer[539]),
      .y(Y[1095]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_321 for neuron1096_1
  function_321 neuron1096_1 (
      .a(~input_layer[2085]),
      .b(input_layer[527]),
      .c(~input_layer[1303]),
      .d(input_layer[269]),
      .e(~input_layer[634]),
      .f(input_layer[1475]),
      .y(Y[1096]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1097_1
  function_64 neuron1097_1 (
      .a(input_layer[2136]),
      .b(input_layer[313]),
      .c(input_layer[1950]),
      .d(~input_layer[994]),
      .e(input_layer[1982]),
      .y(Y[1097]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1098_1
  function_35 neuron1098_1 (
      .a(~input_layer[1503]),
      .b(~input_layer[1456]),
      .c(input_layer[970]),
      .d(~input_layer[1964]),
      .e(input_layer[1852]),
      .y(Y[1098]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1099_1
  function_67 neuron1099_1 (
      .a(input_layer[976]),
      .b(input_layer[2080]),
      .c(~input_layer[1245]),
      .d(~input_layer[1066]),
      .e(~input_layer[804]),
      .y(Y[1099]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1100_1
  function_3 neuron1100_1 (
      .a(input_layer[1041]),
      .b(input_layer[238]),
      .c(~input_layer[1215]),
      .d(input_layer[331]),
      .e(input_layer[508]),
      .y(Y[1100]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1101_1
  function_92 neuron1101_1 (
      .a(input_layer[1584]),
      .b(input_layer[2092]),
      .c(~input_layer[2304]),
      .d(~input_layer[1097]),
      .y(Y[1101]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1102] = 1'b0;

  // instantiate function_322 for neuron1103_1
  function_322 neuron1103_1 (
      .a(input_layer[1381]),
      .b(input_layer[2138]),
      .c(~input_layer[1078]),
      .d(input_layer[696]),
      .e(input_layer[1010]),
      .f(input_layer[394]),
      .y(Y[1103]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1104_1
  function_125 neuron1104_1 (
      .a(~input_layer[2127]),
      .b(~input_layer[1939]),
      .c(input_layer[979]),
      .d(~input_layer[2086]),
      .e(~input_layer[1960]),
      .y(Y[1104]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_123 for neuron1105_1
  function_123 neuron1105_1 (
      .a(~input_layer[478]),
      .b(~input_layer[1456]),
      .c(~input_layer[1380]),
      .d(input_layer[603]),
      .e(input_layer[1562]),
      .f(~input_layer[855]),
      .y(Y[1105]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron1106_1
  function_33 neuron1106_1 (
      .a(~input_layer[1783]),
      .b(~input_layer[1024]),
      .c(~input_layer[894]),
      .d(~input_layer[353]),
      .e(input_layer[488]),
      .y(Y[1106]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron1107_1
  function_156 neuron1107_1 (
      .a(input_layer[1826]),
      .b(~input_layer[472]),
      .c(~input_layer[566]),
      .d(~input_layer[1518]),
      .e(~input_layer[1821]),
      .y(Y[1107]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1108_1
  function_72 neuron1108_1 (
      .a(~input_layer[2052]),
      .b(input_layer[1777]),
      .c(input_layer[1919]),
      .d(~input_layer[103]),
      .e(input_layer[458]),
      .y(Y[1108]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_224 for neuron1109_1
  function_224 neuron1109_1 (
      .a(~input_layer[2120]),
      .b(input_layer[1784]),
      .c(~input_layer[2202]),
      .d(input_layer[1627]),
      .y(Y[1109]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron1110_1
  function_33 neuron1110_1 (
      .a(input_layer[636]),
      .b(input_layer[730]),
      .c(~input_layer[2296]),
      .d(~input_layer[1288]),
      .e(~input_layer[1169]),
      .y(Y[1110]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron1111_1
  function_202 neuron1111_1 (
      .a(input_layer[1134]),
      .b(~input_layer[389]),
      .c(~input_layer[1800]),
      .d(~input_layer[1326]),
      .e(input_layer[1998]),
      .y(Y[1111]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1112_1
  function_139 neuron1112_1 (
      .a(input_layer[1687]),
      .b(~input_layer[649]),
      .c(input_layer[2251]),
      .d(input_layer[1566]),
      .e(~input_layer[1742]),
      .y(Y[1112]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_68 for neuron1113_1
  function_68 neuron1113_1 (
      .a(input_layer[232]),
      .b(~input_layer[1143]),
      .c(~input_layer[1186]),
      .d(~input_layer[1403]),
      .e(~input_layer[900]),
      .f(~input_layer[262]),
      .y(Y[1113]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_323 for neuron1114_1
  function_323 neuron1114_1 (
      .a(~input_layer[1456]),
      .b(input_layer[2113]),
      .c(input_layer[2114]),
      .d(input_layer[1698]),
      .e(~input_layer[2335]),
      .f(input_layer[1938]),
      .y(Y[1114]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1115_1
  function_10 neuron1115_1 (
      .a(input_layer[201]),
      .b(input_layer[1165]),
      .c(~input_layer[614]),
      .d(~input_layer[363]),
      .y(Y[1115]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_324 for neuron1116_1
  function_324 neuron1116_1 (
      .a(input_layer[549]),
      .b(input_layer[1401]),
      .c(input_layer[1869]),
      .d(input_layer[1002]),
      .e(~input_layer[802]),
      .f(input_layer[387]),
      .y(Y[1116]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1117_1
  function_99 neuron1117_1 (
      .a(input_layer[561]),
      .b(input_layer[1862]),
      .c(input_layer[2226]),
      .d(~input_layer[1480]),
      .e(~input_layer[1290]),
      .f(input_layer[1995]),
      .y(Y[1117]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1118_1
  function_307 neuron1118_1 (
      .a(~input_layer[825]),
      .b(~input_layer[582]),
      .c(input_layer[1756]),
      .d(~input_layer[1321]),
      .e(input_layer[185]),
      .y(Y[1118]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1119_1
  function_21 neuron1119_1 (
      .a(~input_layer[994]),
      .b(~input_layer[785]),
      .c(~input_layer[860]),
      .d(input_layer[1131]),
      .y(Y[1119]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1120_1
  function_24 neuron1120_1 (
      .a(~input_layer[1160]),
      .y(Y[1120]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_325 for neuron1121_1
  function_325 neuron1121_1 (
      .a(input_layer[207]),
      .b(~input_layer[699]),
      .c(input_layer[356]),
      .d(input_layer[371]),
      .e(input_layer[915]),
      .f(input_layer[1346]),
      .y(Y[1121]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_198 for neuron1122_1
  function_198 neuron1122_1 (
      .a(~input_layer[1531]),
      .b(input_layer[608]),
      .c(input_layer[1015]),
      .d(~input_layer[1378]),
      .e(input_layer[2329]),
      .y(Y[1122]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1123_1
  function_90 neuron1123_1 (
      .a(~input_layer[1249]),
      .b(input_layer[1836]),
      .c(~input_layer[730]),
      .d(~input_layer[211]),
      .e(~input_layer[1006]),
      .y(Y[1123]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1124_1
  function_18 neuron1124_1 (
      .a(~input_layer[1124]),
      .b(~input_layer[1835]),
      .c(~input_layer[2221]),
      .d(~input_layer[2161]),
      .e(~input_layer[1627]),
      .y(Y[1124]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron1125_1
  function_34 neuron1125_1 (
      .a(input_layer[934]),
      .b(input_layer[2305]),
      .c(input_layer[1358]),
      .d(input_layer[815]),
      .e(~input_layer[922]),
      .y(Y[1125]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_283 for neuron1126_1
  function_283 neuron1126_1 (
      .a(~input_layer[1466]),
      .b(input_layer[693]),
      .c(~input_layer[1595]),
      .d(input_layer[966]),
      .e(~input_layer[1298]),
      .f(input_layer[14]),
      .y(Y[1126]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1127_1
  function_126 neuron1127_1 (
      .a(input_layer[1957]),
      .b(input_layer[1588]),
      .c(~input_layer[1127]),
      .d(~input_layer[204]),
      .e(~input_layer[1404]),
      .y(Y[1127]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1128_1
  function_16 neuron1128_1 (
      .a(input_layer[1526]),
      .b(input_layer[2235]),
      .c(input_layer[535]),
      .y(Y[1128]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1129_1
  function_1 neuron1129_1 (
      .a(~input_layer[1229]),
      .b(~input_layer[233]),
      .c(~input_layer[1376]),
      .d(~input_layer[2024]),
      .e(~input_layer[1567]),
      .f(input_layer[133]),
      .y(Y[1129]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1130_1
  function_54 neuron1130_1 (
      .a(input_layer[373]),
      .b(input_layer[2201]),
      .c(~input_layer[1310]),
      .d(input_layer[594]),
      .e(input_layer[466]),
      .f(~input_layer[1995]),
      .y(Y[1130]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_284 for neuron1131_1
  function_284 neuron1131_1 (
      .a(~input_layer[2312]),
      .b(input_layer[1444]),
      .c(input_layer[1901]),
      .d(input_layer[1504]),
      .e(~input_layer[1526]),
      .f(input_layer[1407]),
      .y(Y[1131]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1132_1
  function_12 neuron1132_1 (
      .a(~input_layer[890]),
      .b(~input_layer[408]),
      .c(~input_layer[513]),
      .y(Y[1132]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1133_1
  function_100 neuron1133_1 (
      .a(input_layer[1034]),
      .b(~input_layer[450]),
      .c(~input_layer[784]),
      .y(Y[1133]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_224 for neuron1134_1
  function_224 neuron1134_1 (
      .a(~input_layer[128]),
      .b(~input_layer[1135]),
      .c(input_layer[2226]),
      .d(~input_layer[2052]),
      .y(Y[1134]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_326 for neuron1135_1
  function_326 neuron1135_1 (
      .a(input_layer[732]),
      .b(~input_layer[411]),
      .c(input_layer[351]),
      .d(input_layer[2334]),
      .e(input_layer[1942]),
      .f(input_layer[887]),
      .y(Y[1135]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1136_1
  function_12 neuron1136_1 (
      .a(~input_layer[1619]),
      .b(~input_layer[825]),
      .c(input_layer[721]),
      .y(Y[1136]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1137_1
  function_63 neuron1137_1 (
      .a(input_layer[1250]),
      .b(~input_layer[885]),
      .c(input_layer[373]),
      .d(input_layer[352]),
      .y(Y[1137]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1138_1
  function_169 neuron1138_1 (
      .a(~input_layer[1410]),
      .b(input_layer[630]),
      .c(input_layer[1503]),
      .d(input_layer[1519]),
      .e(~input_layer[377]),
      .f(~input_layer[428]),
      .y(Y[1138]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1139_1
  function_21 neuron1139_1 (
      .a(~input_layer[607]),
      .b(~input_layer[2158]),
      .c(~input_layer[1351]),
      .d(~input_layer[292]),
      .y(Y[1139]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_327 for neuron1140_1
  function_327 neuron1140_1 (
      .a(~input_layer[737]),
      .b(~input_layer[992]),
      .c(input_layer[1652]),
      .d(input_layer[1431]),
      .e(input_layer[1514]),
      .f(~input_layer[106]),
      .y(Y[1140]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1141_1
  function_25 neuron1141_1 (
      .a(input_layer[2168]),
      .b(input_layer[1250]),
      .c(input_layer[2310]),
      .d(input_layer[1927]),
      .e(input_layer[427]),
      .y(Y[1141]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1142_1
  function_24 neuron1142_1 (
      .a(input_layer[1777]),
      .y(Y[1142]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_328 for neuron1143_1
  function_328 neuron1143_1 (
      .a(~input_layer[649]),
      .b(~input_layer[2145]),
      .c(input_layer[353]),
      .d(input_layer[2169]),
      .e(input_layer[1356]),
      .f(input_layer[187]),
      .y(Y[1143]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1144_1
  function_92 neuron1144_1 (
      .a(input_layer[811]),
      .b(~input_layer[209]),
      .c(input_layer[679]),
      .d(~input_layer[108]),
      .y(Y[1144]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_69 for neuron1145_1
  function_69 neuron1145_1 (
      .a(input_layer[892]),
      .b(~input_layer[302]),
      .c(input_layer[932]),
      .d(~input_layer[1249]),
      .e(input_layer[2314]),
      .y(Y[1145]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1146_1
  function_56 neuron1146_1 (
      .a(~input_layer[862]),
      .b(input_layer[688]),
      .c(~input_layer[132]),
      .d(~input_layer[140]),
      .e(input_layer[1650]),
      .y(Y[1146]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1147] = 1'b0;

  // instantiate function_11 for neuron1148_1
  function_11 neuron1148_1 (
      .a(input_layer[1074]),
      .b(~input_layer[1917]),
      .c(input_layer[1364]),
      .d(input_layer[2295]),
      .y(Y[1148]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1149_1
  function_107 neuron1149_1 (
      .a(~input_layer[522]),
      .b(~input_layer[2239]),
      .c(input_layer[1003]),
      .d(~input_layer[1087]),
      .y(Y[1149]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1150_1
  function_16 neuron1150_1 (
      .a(input_layer[2232]),
      .b(input_layer[1382]),
      .c(input_layer[1261]),
      .y(Y[1150]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_111 for neuron1151_1
  function_111 neuron1151_1 (
      .a(input_layer[1982]),
      .b(~input_layer[1751]),
      .c(~input_layer[1663]),
      .d(input_layer[1726]),
      .e(~input_layer[2294]),
      .f(~input_layer[205]),
      .y(Y[1151]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1152_1
  function_25 neuron1152_1 (
      .a(input_layer[407]),
      .b(input_layer[519]),
      .c(input_layer[189]),
      .d(input_layer[578]),
      .e(~input_layer[451]),
      .y(Y[1152]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1153_1
  function_162 neuron1153_1 (
      .a(~input_layer[1782]),
      .b(~input_layer[2037]),
      .c(~input_layer[1772]),
      .d(~input_layer[1329]),
      .e(input_layer[888]),
      .y(Y[1153]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1154_1
  function_5 neuron1154_1 (
      .a(input_layer[1542]),
      .b(input_layer[1465]),
      .y(Y[1154]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1155_1
  function_169 neuron1155_1 (
      .a(input_layer[2223]),
      .b(~input_layer[1456]),
      .c(input_layer[2051]),
      .d(~input_layer[905]),
      .e(input_layer[856]),
      .f(input_layer[1719]),
      .y(Y[1155]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_172 for neuron1156_1
  function_172 neuron1156_1 (
      .a(~input_layer[771]),
      .b(input_layer[956]),
      .c(~input_layer[131]),
      .d(input_layer[96]),
      .e(~input_layer[932]),
      .f(input_layer[1712]),
      .y(Y[1156]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1157_1
  function_12 neuron1157_1 (
      .a(~input_layer[951]),
      .b(~input_layer[1900]),
      .c(~input_layer[627]),
      .y(Y[1157]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1158_1
  function_11 neuron1158_1 (
      .a(input_layer[307]),
      .b(input_layer[283]),
      .c(input_layer[1769]),
      .d(~input_layer[1969]),
      .y(Y[1158]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1159_1
  function_116 neuron1159_1 (
      .a(input_layer[1705]),
      .b(input_layer[2061]),
      .c(input_layer[2162]),
      .d(input_layer[1305]),
      .y(Y[1159]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1160_1
  function_104 neuron1160_1 (
      .a(input_layer[2207]),
      .b(~input_layer[1701]),
      .c(~input_layer[1589]),
      .y(Y[1160]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_329 for neuron1161_1
  function_329 neuron1161_1 (
      .a(input_layer[1138]),
      .b(~input_layer[1485]),
      .c(~input_layer[1231]),
      .d(~input_layer[142]),
      .e(input_layer[2096]),
      .f(~input_layer[154]),
      .y(Y[1161]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1162_1
  function_25 neuron1162_1 (
      .a(input_layer[869]),
      .b(input_layer[1821]),
      .c(input_layer[2229]),
      .d(input_layer[682]),
      .e(input_layer[151]),
      .y(Y[1162]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1163_1
  function_146 neuron1163_1 (
      .a(input_layer[454]),
      .b(~input_layer[799]),
      .c(input_layer[1770]),
      .d(~input_layer[851]),
      .e(input_layer[1431]),
      .y(Y[1163]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1164_1
  function_154 neuron1164_1 (
      .a(input_layer[849]),
      .b(~input_layer[1748]),
      .c(input_layer[940]),
      .d(~input_layer[1733]),
      .e(input_layer[2314]),
      .y(Y[1164]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_247 for neuron1165_1
  function_247 neuron1165_1 (
      .a(~input_layer[569]),
      .b(input_layer[2295]),
      .c(~input_layer[777]),
      .d(~input_layer[1786]),
      .e(input_layer[1410]),
      .y(Y[1165]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1166_1
  function_330 neuron1166_1 (
      .a(input_layer[686]),
      .b(input_layer[1182]),
      .c(input_layer[1148]),
      .d(input_layer[596]),
      .e(~input_layer[995]),
      .f(input_layer[155]),
      .y(Y[1166]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1167_1
  function_154 neuron1167_1 (
      .a(input_layer[1492]),
      .b(input_layer[1413]),
      .c(~input_layer[607]),
      .d(~input_layer[793]),
      .e(~input_layer[685]),
      .y(Y[1167]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1168_1
  function_139 neuron1168_1 (
      .a(input_layer[1461]),
      .b(input_layer[2065]),
      .c(input_layer[1909]),
      .d(~input_layer[1734]),
      .e(~input_layer[844]),
      .y(Y[1168]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1169_1
  function_5 neuron1169_1 (
      .a(input_layer[902]),
      .b(input_layer[1634]),
      .y(Y[1169]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1170_1
  function_5 neuron1170_1 (
      .a(~input_layer[541]),
      .b(input_layer[226]),
      .y(Y[1170]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1171_1
  function_4 neuron1171_1 (
      .a(input_layer[521]),
      .b(~input_layer[800]),
      .c(input_layer[1956]),
      .d(~input_layer[792]),
      .e(input_layer[802]),
      .y(Y[1171]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1172_1
  function_307 neuron1172_1 (
      .a(~input_layer[411]),
      .b(input_layer[1614]),
      .c(input_layer[2044]),
      .d(input_layer[2140]),
      .e(~input_layer[2257]),
      .y(Y[1172]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_75 for neuron1173_1
  function_75 neuron1173_1 (
      .a(~input_layer[1109]),
      .b(input_layer[1947]),
      .c(input_layer[1941]),
      .d(~input_layer[1120]),
      .e(~input_layer[2007]),
      .y(Y[1173]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1174_1
  function_107 neuron1174_1 (
      .a(~input_layer[450]),
      .b(~input_layer[212]),
      .c(input_layer[1293]),
      .d(~input_layer[824]),
      .y(Y[1174]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1175_1
  function_44 neuron1175_1 (
      .a(~input_layer[2308]),
      .b(input_layer[114]),
      .c(~input_layer[2229]),
      .y(Y[1175]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_331 for neuron1176_1
  function_331 neuron1176_1 (
      .a(~input_layer[811]),
      .b(input_layer[1938]),
      .c(~input_layer[743]),
      .d(input_layer[837]),
      .e(input_layer[153]),
      .y(Y[1176]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1177_1
  function_116 neuron1177_1 (
      .a(input_layer[461]),
      .b(input_layer[650]),
      .c(input_layer[761]),
      .d(~input_layer[531]),
      .y(Y[1177]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_77 for neuron1178_1
  function_77 neuron1178_1 (
      .a(input_layer[1043]),
      .b(~input_layer[2311]),
      .c(input_layer[559]),
      .d(input_layer[1686]),
      .e(input_layer[1601]),
      .f(~input_layer[837]),
      .y(Y[1178]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1179_1
  function_16 neuron1179_1 (
      .a(input_layer[206]),
      .b(~input_layer[827]),
      .c(input_layer[210]),
      .y(Y[1179]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1180_1
  function_18 neuron1180_1 (
      .a(~input_layer[1881]),
      .b(~input_layer[200]),
      .c(~input_layer[1096]),
      .d(~input_layer[2328]),
      .e(~input_layer[2293]),
      .y(Y[1180]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1181_1
  function_54 neuron1181_1 (
      .a(input_layer[2062]),
      .b(input_layer[2031]),
      .c(input_layer[224]),
      .d(~input_layer[1464]),
      .e(input_layer[907]),
      .f(input_layer[2337]),
      .y(Y[1181]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron1182_1
  function_117 neuron1182_1 (
      .a(~input_layer[1142]),
      .b(~input_layer[665]),
      .c(input_layer[1334]),
      .d(~input_layer[1062]),
      .e(~input_layer[1686]),
      .f(~input_layer[2198]),
      .y(Y[1182]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron1183_1
  function_234 neuron1183_1 (
      .a(~input_layer[1688]),
      .b(~input_layer[2113]),
      .c(input_layer[1904]),
      .d(input_layer[561]),
      .e(~input_layer[1679]),
      .f(~input_layer[1628]),
      .y(Y[1183]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1184_1
  function_5 neuron1184_1 (
      .a(~input_layer[541]),
      .b(input_layer[946]),
      .y(Y[1184]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1185_1
  function_11 neuron1185_1 (
      .a(input_layer[828]),
      .b(input_layer[2038]),
      .c(input_layer[1088]),
      .d(input_layer[1575]),
      .y(Y[1185]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1186_1
  function_319 neuron1186_1 (
      .a(input_layer[1303]),
      .b(input_layer[2200]),
      .c(input_layer[1096]),
      .d(input_layer[1280]),
      .e(~input_layer[821]),
      .f(input_layer[297]),
      .y(Y[1186]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1187_1
  function_4 neuron1187_1 (
      .a(input_layer[653]),
      .b(~input_layer[1329]),
      .c(input_layer[267]),
      .d(~input_layer[1332]),
      .e(input_layer[1164]),
      .y(Y[1187]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_160 for neuron1188_1
  function_160 neuron1188_1 (
      .a(input_layer[579]),
      .b(~input_layer[392]),
      .c(input_layer[2242]),
      .d(~input_layer[378]),
      .e(~input_layer[447]),
      .y(Y[1188]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_241 for neuron1189_1
  function_241 neuron1189_1 (
      .a(~input_layer[1282]),
      .b(~input_layer[1188]),
      .c(input_layer[750]),
      .d(~input_layer[2319]),
      .e(input_layer[344]),
      .f(input_layer[1720]),
      .y(Y[1189]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_332 for neuron1190_1
  function_332 neuron1190_1 (
      .a(~input_layer[1630]),
      .b(input_layer[1054]),
      .c(~input_layer[375]),
      .d(~input_layer[774]),
      .e(~input_layer[268]),
      .f(input_layer[2051]),
      .y(Y[1190]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1191_1
  function_12 neuron1191_1 (
      .a(~input_layer[700]),
      .b(~input_layer[225]),
      .c(~input_layer[748]),
      .y(Y[1191]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron1192_1
  function_248 neuron1192_1 (
      .a(~input_layer[1128]),
      .b(~input_layer[1327]),
      .c(~input_layer[410]),
      .d(~input_layer[1238]),
      .e(input_layer[188]),
      .f(input_layer[1182]),
      .y(Y[1192]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_333 for neuron1193_1
  function_333 neuron1193_1 (
      .a(~input_layer[1543]),
      .b(input_layer[1114]),
      .c(input_layer[2025]),
      .d(input_layer[1258]),
      .e(~input_layer[264]),
      .f(~input_layer[1335]),
      .y(Y[1193]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1194_1
  function_44 neuron1194_1 (
      .a(~input_layer[1280]),
      .b(input_layer[1405]),
      .c(input_layer[1854]),
      .y(Y[1194]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1195_1
  function_334 neuron1195_1 (
      .a(~input_layer[665]),
      .b(input_layer[1870]),
      .c(input_layer[963]),
      .d(input_layer[1525]),
      .e(input_layer[1875]),
      .f(input_layer[1410]),
      .y(Y[1195]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1196_1
  function_90 neuron1196_1 (
      .a(~input_layer[1467]),
      .b(input_layer[1960]),
      .c(input_layer[656]),
      .d(~input_layer[1235]),
      .e(~input_layer[262]),
      .y(Y[1196]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1197_1
  function_3 neuron1197_1 (
      .a(input_layer[444]),
      .b(input_layer[429]),
      .c(input_layer[1824]),
      .d(input_layer[330]),
      .e(input_layer[1816]),
      .y(Y[1197]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_160 for neuron1198_1
  function_160 neuron1198_1 (
      .a(input_layer[2324]),
      .b(~input_layer[1283]),
      .c(~input_layer[2146]),
      .d(~input_layer[302]),
      .e(input_layer[2059]),
      .y(Y[1198]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_335 for neuron1199_1
  function_335 neuron1199_1 (
      .a(input_layer[1760]),
      .b(input_layer[1890]),
      .c(input_layer[1279]),
      .d(input_layer[646]),
      .e(input_layer[418]),
      .f(input_layer[2189]),
      .y(Y[1199]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1200_1
  function_18 neuron1200_1 (
      .a(~input_layer[956]),
      .b(~input_layer[1388]),
      .c(~input_layer[286]),
      .d(input_layer[1209]),
      .e(~input_layer[2111]),
      .y(Y[1200]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_336 for neuron1201_1
  function_336 neuron1201_1 (
      .a(input_layer[1588]),
      .b(input_layer[1798]),
      .c(input_layer[1283]),
      .d(~input_layer[2154]),
      .e(~input_layer[638]),
      .f(input_layer[1643]),
      .y(Y[1201]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1202_1
  function_19 neuron1202_1 (
      .a(~input_layer[2130]),
      .b(input_layer[1959]),
      .c(input_layer[208]),
      .d(input_layer[100]),
      .y(Y[1202]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1203_1
  function_14 neuron1203_1 (
      .a(~input_layer[829]),
      .b(~input_layer[2068]),
      .c(~input_layer[1772]),
      .d(input_layer[1536]),
      .e(input_layer[1461]),
      .y(Y[1203]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1204_1
  function_148 neuron1204_1 (
      .a(~input_layer[201]),
      .b(input_layer[537]),
      .c(~input_layer[111]),
      .d(input_layer[896]),
      .y(Y[1204]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1205_1
  function_25 neuron1205_1 (
      .a(input_layer[387]),
      .b(input_layer[393]),
      .c(input_layer[439]),
      .d(input_layer[224]),
      .e(input_layer[413]),
      .y(Y[1205]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1206_1
  function_24 neuron1206_1 (
      .a(input_layer[1193]),
      .y(Y[1206]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_199 for neuron1207_1
  function_199 neuron1207_1 (
      .a(~input_layer[1123]),
      .b(input_layer[2305]),
      .c(~input_layer[1036]),
      .d(~input_layer[205]),
      .e(input_layer[1719]),
      .f(input_layer[1466]),
      .y(Y[1207]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1208_1
  function_3 neuron1208_1 (
      .a(input_layer[1389]),
      .b(input_layer[1307]),
      .c(input_layer[315]),
      .d(input_layer[307]),
      .e(~input_layer[653]),
      .y(Y[1208]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_337 for neuron1209_1
  function_337 neuron1209_1 (
      .a(~input_layer[668]),
      .b(input_layer[1365]),
      .c(~input_layer[404]),
      .d(~input_layer[1402]),
      .e(~input_layer[2193]),
      .f(~input_layer[710]),
      .y(Y[1209]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1210_1
  function_18 neuron1210_1 (
      .a(~input_layer[979]),
      .b(~input_layer[2143]),
      .c(~input_layer[318]),
      .d(~input_layer[1073]),
      .e(~input_layer[354]),
      .y(Y[1210]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1211_1
  function_63 neuron1211_1 (
      .a(input_layer[292]),
      .b(~input_layer[1077]),
      .c(input_layer[941]),
      .d(input_layer[1357]),
      .y(Y[1211]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1212_1
  function_11 neuron1212_1 (
      .a(input_layer[2160]),
      .b(input_layer[1184]),
      .c(input_layer[1506]),
      .d(~input_layer[1916]),
      .y(Y[1212]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1213_1
  function_11 neuron1213_1 (
      .a(input_layer[1827]),
      .b(input_layer[1003]),
      .c(input_layer[1438]),
      .d(input_layer[1641]),
      .y(Y[1213]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron1214_1
  function_152 neuron1214_1 (
      .a(~input_layer[525]),
      .b(input_layer[1918]),
      .c(~input_layer[392]),
      .d(input_layer[2138]),
      .e(~input_layer[902]),
      .f(input_layer[1897]),
      .y(Y[1214]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1215_1
  function_3 neuron1215_1 (
      .a(input_layer[1827]),
      .b(input_layer[1666]),
      .c(input_layer[528]),
      .d(input_layer[867]),
      .e(input_layer[1442]),
      .y(Y[1215]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1216_1
  function_63 neuron1216_1 (
      .a(input_layer[205]),
      .b(input_layer[459]),
      .c(input_layer[1090]),
      .d(input_layer[1388]),
      .y(Y[1216]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_255 for neuron1217_1
  function_255 neuron1217_1 (
      .a(~input_layer[1647]),
      .b(input_layer[2082]),
      .c(input_layer[992]),
      .d(input_layer[393]),
      .e(input_layer[1801]),
      .y(Y[1217]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1218_1
  function_44 neuron1218_1 (
      .a(~input_layer[1253]),
      .b(~input_layer[1789]),
      .c(~input_layer[1454]),
      .y(Y[1218]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1219_1
  function_18 neuron1219_1 (
      .a(~input_layer[769]),
      .b(~input_layer[849]),
      .c(input_layer[2224]),
      .d(~input_layer[279]),
      .e(~input_layer[1171]),
      .y(Y[1219]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1220_1
  function_12 neuron1220_1 (
      .a(~input_layer[1987]),
      .b(~input_layer[1208]),
      .c(~input_layer[210]),
      .y(Y[1220]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1221_1
  function_18 neuron1221_1 (
      .a(~input_layer[815]),
      .b(~input_layer[1700]),
      .c(~input_layer[1580]),
      .d(~input_layer[1167]),
      .e(~input_layer[308]),
      .y(Y[1221]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1222_1
  function_16 neuron1222_1 (
      .a(input_layer[1277]),
      .b(input_layer[486]),
      .c(~input_layer[625]),
      .y(Y[1222]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1223_1
  function_125 neuron1223_1 (
      .a(~input_layer[1694]),
      .b(~input_layer[2314]),
      .c(~input_layer[670]),
      .d(input_layer[1191]),
      .e(input_layer[1166]),
      .y(Y[1223]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_338 for neuron1224_1
  function_338 neuron1224_1 (
      .a(~input_layer[608]),
      .b(input_layer[877]),
      .c(input_layer[2288]),
      .d(input_layer[1575]),
      .e(~input_layer[2130]),
      .f(~input_layer[1399]),
      .y(Y[1224]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1225_1
  function_10 neuron1225_1 (
      .a(input_layer[852]),
      .b(input_layer[2305]),
      .c(input_layer[782]),
      .d(~input_layer[1073]),
      .y(Y[1225]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_339 for neuron1226_1
  function_339 neuron1226_1 (
      .a(~input_layer[1946]),
      .b(~input_layer[1654]),
      .c(input_layer[742]),
      .d(input_layer[835]),
      .e(input_layer[1124]),
      .f(~input_layer[1181]),
      .y(Y[1226]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_122 for neuron1227_1
  function_122 neuron1227_1 (
      .a(~input_layer[438]),
      .b(input_layer[409]),
      .c(~input_layer[1560]),
      .d(input_layer[1008]),
      .e(~input_layer[727]),
      .f(~input_layer[1870]),
      .y(Y[1227]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron1228_1
  function_133 neuron1228_1 (
      .a(~input_layer[831]),
      .b(input_layer[895]),
      .c(input_layer[1014]),
      .d(input_layer[1635]),
      .e(input_layer[297]),
      .y(Y[1228]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_329 for neuron1229_1
  function_329 neuron1229_1 (
      .a(~input_layer[970]),
      .b(input_layer[1120]),
      .c(~input_layer[611]),
      .d(~input_layer[2200]),
      .e(~input_layer[1311]),
      .f(~input_layer[2315]),
      .y(Y[1229]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_266 for neuron1230_1
  function_266 neuron1230_1 (
      .a(~input_layer[319]),
      .b(~input_layer[959]),
      .c(~input_layer[2053]),
      .d(~input_layer[1210]),
      .e(input_layer[1067]),
      .f(~input_layer[306]),
      .y(Y[1230]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_128 for neuron1231_1
  function_128 neuron1231_1 (
      .a(input_layer[1026]),
      .b(~input_layer[1827]),
      .c(~input_layer[2023]),
      .d(input_layer[125]),
      .y(Y[1231]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1232_1
  function_44 neuron1232_1 (
      .a(~input_layer[2240]),
      .b(input_layer[874]),
      .c(input_layer[1418]),
      .y(Y[1232]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1233_1
  function_91 neuron1233_1 (
      .a(input_layer[2034]),
      .b(input_layer[1456]),
      .c(input_layer[1011]),
      .d(input_layer[1346]),
      .e(input_layer[1009]),
      .f(~input_layer[1765]),
      .y(Y[1233]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1234_1
  function_113 neuron1234_1 (
      .a(input_layer[1441]),
      .b(input_layer[617]),
      .c(~input_layer[1558]),
      .d(input_layer[1643]),
      .e(input_layer[880]),
      .f(input_layer[2096]),
      .y(Y[1234]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_287 for neuron1235_1
  function_287 neuron1235_1 (
      .a(~input_layer[2122]),
      .b(~input_layer[1950]),
      .c(~input_layer[2252]),
      .d(input_layer[1891]),
      .e(~input_layer[1829]),
      .f(input_layer[626]),
      .y(Y[1235]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_221 for neuron1236_1
  function_221 neuron1236_1 (
      .a(input_layer[456]),
      .b(~input_layer[1184]),
      .c(~input_layer[1726]),
      .d(~input_layer[295]),
      .e(input_layer[517]),
      .f(input_layer[51]),
      .y(Y[1236]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1237_1
  function_107 neuron1237_1 (
      .a(~input_layer[1800]),
      .b(~input_layer[1256]),
      .c(~input_layer[1412]),
      .d(input_layer[1104]),
      .y(Y[1237]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1238_1
  function_76 neuron1238_1 (
      .a(~input_layer[2134]),
      .b(~input_layer[736]),
      .c(~input_layer[1996]),
      .d(input_layer[1639]),
      .e(~input_layer[1980]),
      .f(~input_layer[1805]),
      .y(Y[1238]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_340 for neuron1239_1
  function_340 neuron1239_1 (
      .a(~input_layer[1103]),
      .b(~input_layer[1122]),
      .c(input_layer[778]),
      .d(input_layer[779]),
      .e(~input_layer[1092]),
      .f(~input_layer[30]),
      .y(Y[1239]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1240_1
  function_12 neuron1240_1 (
      .a(~input_layer[951]),
      .b(~input_layer[2080]),
      .c(~input_layer[2235]),
      .y(Y[1240]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_318 for neuron1241_1
  function_318 neuron1241_1 (
      .a(~input_layer[574]),
      .b(input_layer[1579]),
      .c(input_layer[1140]),
      .d(input_layer[140]),
      .e(~input_layer[655]),
      .f(input_layer[472]),
      .y(Y[1241]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1242_1
  function_11 neuron1242_1 (
      .a(input_layer[1747]),
      .b(input_layer[453]),
      .c(~input_layer[689]),
      .d(input_layer[461]),
      .y(Y[1242]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron1243_1
  function_62 neuron1243_1 (
      .a(input_layer[1153]),
      .b(input_layer[613]),
      .c(~input_layer[2009]),
      .d(~input_layer[704]),
      .y(Y[1243]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1244_1
  function_146 neuron1244_1 (
      .a(input_layer[2032]),
      .b(input_layer[803]),
      .c(input_layer[2317]),
      .d(~input_layer[1834]),
      .e(input_layer[452]),
      .y(Y[1244]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1245_1
  function_10 neuron1245_1 (
      .a(input_layer[1522]),
      .b(input_layer[2161]),
      .c(~input_layer[1283]),
      .d(input_layer[1582]),
      .y(Y[1245]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1246_1
  function_116 neuron1246_1 (
      .a(input_layer[1751]),
      .b(~input_layer[780]),
      .c(input_layer[1256]),
      .d(input_layer[1441]),
      .y(Y[1246]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1247_1
  function_45 neuron1247_1 (
      .a(~input_layer[1414]),
      .b(~input_layer[448]),
      .c(~input_layer[1527]),
      .d(~input_layer[1059]),
      .e(~input_layer[2305]),
      .f(~input_layer[1899]),
      .y(Y[1247]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1248_1
  function_12 neuron1248_1 (
      .a(~input_layer[1191]),
      .b(~input_layer[192]),
      .c(~input_layer[1311]),
      .y(Y[1248]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_341 for neuron1249_1
  function_341 neuron1249_1 (
      .a(input_layer[2229]),
      .b(input_layer[120]),
      .c(~input_layer[955]),
      .d(~input_layer[1193]),
      .e(input_layer[1814]),
      .f(input_layer[261]),
      .y(Y[1249]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1250_1
  function_37 neuron1250_1 (
      .a(input_layer[744]),
      .b(input_layer[1548]),
      .c(~input_layer[292]),
      .d(~input_layer[813]),
      .e(input_layer[2012]),
      .y(Y[1250]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1251_1
  function_67 neuron1251_1 (
      .a(input_layer[547]),
      .b(input_layer[661]),
      .c(input_layer[2092]),
      .d(~input_layer[2145]),
      .e(~input_layer[949]),
      .y(Y[1251]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_207 for neuron1252_1
  function_207 neuron1252_1 (
      .a(~input_layer[636]),
      .b(input_layer[904]),
      .c(input_layer[1959]),
      .d(~input_layer[1105]),
      .e(~input_layer[960]),
      .f(~input_layer[1700]),
      .y(Y[1252]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1253_1
  function_40 neuron1253_1 (
      .a(~input_layer[484]),
      .b(~input_layer[1716]),
      .c(~input_layer[354]),
      .d(input_layer[631]),
      .e(~input_layer[223]),
      .f(~input_layer[1086]),
      .y(Y[1253]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1254_1
  function_99 neuron1254_1 (
      .a(input_layer[1003]),
      .b(input_layer[2295]),
      .c(~input_layer[1383]),
      .d(input_layer[1061]),
      .e(input_layer[1277]),
      .f(~input_layer[2178]),
      .y(Y[1254]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1255_1
  function_63 neuron1255_1 (
      .a(input_layer[1552]),
      .b(~input_layer[1613]),
      .c(input_layer[569]),
      .d(input_layer[1260]),
      .y(Y[1255]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1256_1
  function_87 neuron1256_1 (
      .a(input_layer[1245]),
      .b(input_layer[1204]),
      .c(input_layer[1593]),
      .d(~input_layer[1323]),
      .e(input_layer[1308]),
      .f(~input_layer[2133]),
      .y(Y[1256]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1257_1
  function_12 neuron1257_1 (
      .a(~input_layer[2115]),
      .b(~input_layer[305]),
      .c(input_layer[639]),
      .y(Y[1257]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_153 for neuron1258_1
  function_153 neuron1258_1 (
      .a(~input_layer[1965]),
      .b(input_layer[2000]),
      .c(input_layer[1377]),
      .d(input_layer[1349]),
      .e(~input_layer[1332]),
      .f(input_layer[1193]),
      .y(Y[1258]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1259_1
  function_54 neuron1259_1 (
      .a(input_layer[1409]),
      .b(input_layer[1320]),
      .c(input_layer[593]),
      .d(input_layer[1169]),
      .e(input_layer[1525]),
      .f(input_layer[1419]),
      .y(Y[1259]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron1260_1
  function_234 neuron1260_1 (
      .a(input_layer[495]),
      .b(~input_layer[2213]),
      .c(~input_layer[863]),
      .d(~input_layer[1027]),
      .e(~input_layer[1930]),
      .f(~input_layer[1954]),
      .y(Y[1260]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1261_1
  function_319 neuron1261_1 (
      .a(input_layer[870]),
      .b(input_layer[830]),
      .c(input_layer[1747]),
      .d(~input_layer[1903]),
      .e(input_layer[856]),
      .f(input_layer[1716]),
      .y(Y[1261]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1262_1
  function_149 neuron1262_1 (
      .a(~input_layer[1452]),
      .b(~input_layer[1492]),
      .c(~input_layer[329]),
      .d(input_layer[2141]),
      .y(Y[1262]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1263_1
  function_12 neuron1263_1 (
      .a(~input_layer[662]),
      .b(~input_layer[806]),
      .c(~input_layer[119]),
      .y(Y[1263]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_118 for neuron1264_1
  function_118 neuron1264_1 (
      .a(input_layer[1509]),
      .b(input_layer[1119]),
      .c(~input_layer[2293]),
      .d(input_layer[418]),
      .e(input_layer[1139]),
      .y(Y[1264]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1265_1
  function_40 neuron1265_1 (
      .a(~input_layer[550]),
      .b(~input_layer[1590]),
      .c(~input_layer[2324]),
      .d(input_layer[1056]),
      .e(~input_layer[591]),
      .f(~input_layer[1516]),
      .y(Y[1265]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1266_1
  function_116 neuron1266_1 (
      .a(~input_layer[472]),
      .b(input_layer[764]),
      .c(input_layer[2241]),
      .d(input_layer[1242]),
      .y(Y[1266]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1267_1
  function_11 neuron1267_1 (
      .a(input_layer[1418]),
      .b(input_layer[1787]),
      .c(input_layer[678]),
      .d(input_layer[1298]),
      .y(Y[1267]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_342 for neuron1268_1
  function_342 neuron1268_1 (
      .a(input_layer[884]),
      .b(~input_layer[1983]),
      .c(input_layer[1719]),
      .d(~input_layer[577]),
      .e(input_layer[2201]),
      .f(input_layer[2158]),
      .y(Y[1268]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1269_1
  function_16 neuron1269_1 (
      .a(input_layer[1949]),
      .b(input_layer[353]),
      .c(~input_layer[1823]),
      .y(Y[1269]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_343 for neuron1270_1
  function_343 neuron1270_1 (
      .a(~input_layer[907]),
      .b(input_layer[750]),
      .c(input_layer[2078]),
      .d(input_layer[1637]),
      .e(~input_layer[2196]),
      .f(input_layer[2252]),
      .y(Y[1270]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1271_1
  function_26 neuron1271_1 (
      .a(input_layer[1385]),
      .b(~input_layer[993]),
      .y(Y[1271]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1272_1
  function_319 neuron1272_1 (
      .a(input_layer[211]),
      .b(~input_layer[1767]),
      .c(input_layer[183]),
      .d(input_layer[477]),
      .e(input_layer[154]),
      .f(input_layer[188]),
      .y(Y[1272]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_291 for neuron1273_1
  function_291 neuron1273_1 (
      .a(input_layer[1740]),
      .b(~input_layer[2310]),
      .c(~input_layer[2050]),
      .d(input_layer[537]),
      .e(~input_layer[869]),
      .f(input_layer[153]),
      .y(Y[1273]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1274_1
  function_21 neuron1274_1 (
      .a(~input_layer[1374]),
      .b(~input_layer[1250]),
      .c(~input_layer[1190]),
      .d(input_layer[1884]),
      .y(Y[1274]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1275_1
  function_5 neuron1275_1 (
      .a(input_layer[1585]),
      .b(~input_layer[1053]),
      .y(Y[1275]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_124 for neuron1276_1
  function_124 neuron1276_1 (
      .a(~input_layer[1069]),
      .b(input_layer[826]),
      .c(~input_layer[600]),
      .d(input_layer[743]),
      .e(input_layer[1427]),
      .f(input_layer[335]),
      .y(Y[1276]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_344 for neuron1277_1
  function_344 neuron1277_1 (
      .a(input_layer[1101]),
      .b(~input_layer[1732]),
      .c(~input_layer[221]),
      .d(input_layer[2059]),
      .e(input_layer[477]),
      .f(input_layer[465]),
      .y(Y[1277]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1278_1
  function_298 neuron1278_1 (
      .a(input_layer[1243]),
      .b(~input_layer[1704]),
      .c(~input_layer[864]),
      .d(input_layer[1241]),
      .e(~input_layer[1336]),
      .y(Y[1278]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_48 for neuron1279_1
  function_48 neuron1279_1 (
      .a(input_layer[1398]),
      .b(input_layer[1146]),
      .c(~input_layer[617]),
      .d(~input_layer[1580]),
      .e(~input_layer[1260]),
      .y(Y[1279]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron1280_1
  function_132 neuron1280_1 (
      .a(~input_layer[1873]),
      .b(input_layer[1568]),
      .c(input_layer[1736]),
      .d(input_layer[468]),
      .e(~input_layer[1906]),
      .y(Y[1280]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_345 for neuron1281_1
  function_345 neuron1281_1 (
      .a(input_layer[856]),
      .b(~input_layer[1315]),
      .c(input_layer[473]),
      .d(~input_layer[1186]),
      .e(~input_layer[1342]),
      .f(~input_layer[695]),
      .y(Y[1281]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1282_1
  function_162 neuron1282_1 (
      .a(~input_layer[204]),
      .b(~input_layer[1450]),
      .c(input_layer[1301]),
      .d(~input_layer[680]),
      .e(~input_layer[2254]),
      .y(Y[1282]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1283_1
  function_100 neuron1283_1 (
      .a(~input_layer[1627]),
      .b(input_layer[2151]),
      .c(input_layer[794]),
      .y(Y[1283]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1284_1
  function_3 neuron1284_1 (
      .a(input_layer[1486]),
      .b(input_layer[1508]),
      .c(input_layer[1774]),
      .d(input_layer[1897]),
      .e(input_layer[1868]),
      .y(Y[1284]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1285_1
  function_21 neuron1285_1 (
      .a(~input_layer[1802]),
      .b(~input_layer[1673]),
      .c(~input_layer[1702]),
      .d(~input_layer[1701]),
      .y(Y[1285]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1286_1
  function_67 neuron1286_1 (
      .a(~input_layer[808]),
      .b(input_layer[1622]),
      .c(input_layer[1037]),
      .d(input_layer[1330]),
      .e(input_layer[1575]),
      .y(Y[1286]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1287_1
  function_99 neuron1287_1 (
      .a(input_layer[1828]),
      .b(input_layer[1339]),
      .c(~input_layer[1137]),
      .d(input_layer[671]),
      .e(input_layer[37]),
      .f(input_layer[1947]),
      .y(Y[1287]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1288_1
  function_11 neuron1288_1 (
      .a(input_layer[445]),
      .b(input_layer[2121]),
      .c(input_layer[777]),
      .d(~input_layer[1242]),
      .y(Y[1288]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_74 for neuron1289_1
  function_74 neuron1289_1 (
      .a(~input_layer[1366]),
      .b(~input_layer[435]),
      .c(input_layer[1894]),
      .d(input_layer[1825]),
      .e(input_layer[755]),
      .y(Y[1289]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1290_1
  function_116 neuron1290_1 (
      .a(input_layer[2141]),
      .b(input_layer[2210]),
      .c(input_layer[2142]),
      .d(~input_layer[1889]),
      .y(Y[1290]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1291_1
  function_11 neuron1291_1 (
      .a(input_layer[1294]),
      .b(input_layer[1116]),
      .c(input_layer[979]),
      .d(input_layer[976]),
      .y(Y[1291]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_105 for neuron1292_1
  function_105 neuron1292_1 (
      .a(input_layer[813]),
      .b(~input_layer[313]),
      .c(~input_layer[395]),
      .d(~input_layer[196]),
      .e(input_layer[1706]),
      .f(~input_layer[2269]),
      .y(Y[1292]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_141 for neuron1293_1
  function_141 neuron1293_1 (
      .a(input_layer[1198]),
      .b(input_layer[1039]),
      .c(~input_layer[277]),
      .d(~input_layer[544]),
      .e(input_layer[1125]),
      .f(~input_layer[976]),
      .y(Y[1293]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1294_1
  function_162 neuron1294_1 (
      .a(~input_layer[522]),
      .b(~input_layer[1118]),
      .c(~input_layer[410]),
      .d(~input_layer[1203]),
      .e(input_layer[737]),
      .y(Y[1294]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_346 for neuron1295_1
  function_346 neuron1295_1 (
      .a(~input_layer[1715]),
      .b(~input_layer[1614]),
      .c(input_layer[1882]),
      .d(input_layer[133]),
      .e(input_layer[1084]),
      .f(input_layer[1820]),
      .y(Y[1295]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1296_1
  function_139 neuron1296_1 (
      .a(input_layer[746]),
      .b(~input_layer[1523]),
      .c(~input_layer[717]),
      .d(input_layer[2075]),
      .e(input_layer[333]),
      .y(Y[1296]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1297_1
  function_26 neuron1297_1 (
      .a(~input_layer[1661]),
      .b(~input_layer[1735]),
      .y(Y[1297]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1298_1
  function_146 neuron1298_1 (
      .a(input_layer[1788]),
      .b(input_layer[934]),
      .c(input_layer[547]),
      .d(~input_layer[733]),
      .e(input_layer[725]),
      .y(Y[1298]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1299_1
  function_21 neuron1299_1 (
      .a(~input_layer[631]),
      .b(~input_layer[2033]),
      .c(~input_layer[2207]),
      .d(~input_layer[1679]),
      .y(Y[1299]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_347 for neuron1300_1
  function_347 neuron1300_1 (
      .a(~input_layer[855]),
      .b(input_layer[1590]),
      .c(input_layer[1362]),
      .d(~input_layer[2037]),
      .e(input_layer[1851]),
      .f(input_layer[1328]),
      .y(Y[1300]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1301_1
  function_181 neuron1301_1 (
      .a(~input_layer[735]),
      .b(~input_layer[357]),
      .c(~input_layer[665]),
      .d(input_layer[382]),
      .e(~input_layer[953]),
      .f(input_layer[402]),
      .y(Y[1301]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron1302_1
  function_303 neuron1302_1 (
      .a(input_layer[933]),
      .b(input_layer[729]),
      .c(input_layer[519]),
      .d(input_layer[2045]),
      .e(~input_layer[1648]),
      .f(~input_layer[135]),
      .y(Y[1302]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1303_1
  function_10 neuron1303_1 (
      .a(input_layer[293]),
      .b(input_layer[1959]),
      .c(~input_layer[494]),
      .d(input_layer[1542]),
      .y(Y[1303]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_207 for neuron1304_1
  function_207 neuron1304_1 (
      .a(input_layer[1380]),
      .b(~input_layer[1645]),
      .c(input_layer[1492]),
      .d(input_layer[1531]),
      .e(~input_layer[717]),
      .f(~input_layer[1701]),
      .y(Y[1304]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron1305_1
  function_33 neuron1305_1 (
      .a(~input_layer[1911]),
      .b(~input_layer[1843]),
      .c(input_layer[313]),
      .d(~input_layer[725]),
      .e(~input_layer[2083]),
      .y(Y[1305]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1306_1
  function_10 neuron1306_1 (
      .a(input_layer[999]),
      .b(input_layer[230]),
      .c(~input_layer[788]),
      .d(~input_layer[1745]),
      .y(Y[1306]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1307_1
  function_54 neuron1307_1 (
      .a(input_layer[2070]),
      .b(~input_layer[1582]),
      .c(input_layer[1810]),
      .d(input_layer[929]),
      .e(input_layer[1187]),
      .f(input_layer[1702]),
      .y(Y[1307]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1308_1
  function_26 neuron1308_1 (
      .a(input_layer[1909]),
      .b(~input_layer[2162]),
      .y(Y[1308]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_348 for neuron1309_1
  function_348 neuron1309_1 (
      .a(input_layer[2308]),
      .b(~input_layer[2209]),
      .c(input_layer[1360]),
      .d(~input_layer[732]),
      .e(~input_layer[703]),
      .f(input_layer[1262]),
      .y(Y[1309]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1310_1
  function_0 neuron1310_1 (
      .a(input_layer[1411]),
      .b(input_layer[197]),
      .c(input_layer[366]),
      .d(input_layer[1724]),
      .e(input_layer[1647]),
      .y(Y[1310]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_349 for neuron1311_1
  function_349 neuron1311_1 (
      .a(~input_layer[1378]),
      .b(input_layer[1327]),
      .c(input_layer[237]),
      .d(~input_layer[531]),
      .e(~input_layer[1010]),
      .f(input_layer[89]),
      .y(Y[1311]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1312_1
  function_21 neuron1312_1 (
      .a(~input_layer[1109]),
      .b(~input_layer[1061]),
      .c(~input_layer[1427]),
      .d(input_layer[572]),
      .y(Y[1312]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1313_1
  function_87 neuron1313_1 (
      .a(input_layer[2234]),
      .b(~input_layer[1059]),
      .c(input_layer[1751]),
      .d(input_layer[181]),
      .e(input_layer[1097]),
      .f(input_layer[99]),
      .y(Y[1313]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1314_1
  function_334 neuron1314_1 (
      .a(input_layer[1470]),
      .b(~input_layer[1789]),
      .c(~input_layer[1770]),
      .d(input_layer[1318]),
      .e(input_layer[1368]),
      .f(~input_layer[2283]),
      .y(Y[1314]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_350 for neuron1315_1
  function_350 neuron1315_1 (
      .a(input_layer[2228]),
      .b(~input_layer[311]),
      .c(~input_layer[1447]),
      .d(~input_layer[440]),
      .e(~input_layer[437]),
      .y(Y[1315]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1316_1
  function_19 neuron1316_1 (
      .a(input_layer[1807]),
      .b(input_layer[1731]),
      .c(input_layer[1823]),
      .d(input_layer[1121]),
      .y(Y[1316]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron1317_1
  function_165 neuron1317_1 (
      .a(~input_layer[1133]),
      .b(~input_layer[2324]),
      .c(input_layer[1192]),
      .d(~input_layer[2094]),
      .e(input_layer[628]),
      .f(~input_layer[882]),
      .y(Y[1317]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1318_1
  function_3 neuron1318_1 (
      .a(input_layer[312]),
      .b(input_layer[1077]),
      .c(input_layer[911]),
      .d(input_layer[1715]),
      .e(input_layer[1031]),
      .y(Y[1318]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1319_1
  function_91 neuron1319_1 (
      .a(input_layer[1943]),
      .b(input_layer[1456]),
      .c(~input_layer[712]),
      .d(input_layer[1845]),
      .e(~input_layer[2339]),
      .f(input_layer[1936]),
      .y(Y[1319]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_351 for neuron1320_1
  function_351 neuron1320_1 (
      .a(~input_layer[1018]),
      .b(input_layer[1987]),
      .c(input_layer[1137]),
      .d(~input_layer[1830]),
      .e(input_layer[191]),
      .f(~input_layer[1309]),
      .y(Y[1320]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1321_1
  function_53 neuron1321_1 (
      .a(input_layer[1784]),
      .b(input_layer[355]),
      .c(~input_layer[273]),
      .d(~input_layer[1070]),
      .e(input_layer[1093]),
      .y(Y[1321]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1322_1
  function_21 neuron1322_1 (
      .a(~input_layer[1246]),
      .b(~input_layer[1146]),
      .c(~input_layer[1356]),
      .d(~input_layer[1425]),
      .y(Y[1322]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1323_1
  function_162 neuron1323_1 (
      .a(~input_layer[970]),
      .b(~input_layer[2061]),
      .c(~input_layer[1419]),
      .d(input_layer[871]),
      .e(~input_layer[1268]),
      .y(Y[1323]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1324_1
  function_10 neuron1324_1 (
      .a(input_layer[748]),
      .b(~input_layer[1794]),
      .c(input_layer[353]),
      .d(~input_layer[180]),
      .y(Y[1324]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1325_1
  function_18 neuron1325_1 (
      .a(~input_layer[286]),
      .b(~input_layer[1360]),
      .c(~input_layer[858]),
      .d(~input_layer[1112]),
      .e(input_layer[468]),
      .y(Y[1325]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1326_1
  function_26 neuron1326_1 (
      .a(~input_layer[1071]),
      .b(~input_layer[1185]),
      .y(Y[1326]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1327_1
  function_125 neuron1327_1 (
      .a(~input_layer[1046]),
      .b(~input_layer[746]),
      .c(input_layer[737]),
      .d(~input_layer[1075]),
      .e(input_layer[1432]),
      .y(Y[1327]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1328_1
  function_231 neuron1328_1 (
      .a(~input_layer[1060]),
      .b(~input_layer[1436]),
      .c(input_layer[474]),
      .d(~input_layer[2072]),
      .e(input_layer[1613]),
      .f(~input_layer[2337]),
      .y(Y[1328]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1329_1
  function_148 neuron1329_1 (
      .a(~input_layer[1030]),
      .b(~input_layer[573]),
      .c(input_layer[284]),
      .d(~input_layer[2055]),
      .y(Y[1329]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron1330_1
  function_65 neuron1330_1 (
      .a(~input_layer[1792]),
      .b(~input_layer[187]),
      .c(~input_layer[1464]),
      .d(input_layer[1115]),
      .e(~input_layer[2115]),
      .f(~input_layer[154]),
      .y(Y[1330]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1331_1
  function_56 neuron1331_1 (
      .a(~input_layer[1642]),
      .b(~input_layer[1445]),
      .c(input_layer[605]),
      .d(~input_layer[1797]),
      .e(~input_layer[1065]),
      .y(Y[1331]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1332_1
  function_91 neuron1332_1 (
      .a(input_layer[1028]),
      .b(input_layer[577]),
      .c(input_layer[887]),
      .d(input_layer[245]),
      .e(input_layer[1610]),
      .f(~input_layer[358]),
      .y(Y[1332]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1333_1
  function_167 neuron1333_1 (
      .a(~input_layer[771]),
      .b(input_layer[595]),
      .c(~input_layer[907]),
      .d(~input_layer[1797]),
      .e(input_layer[979]),
      .y(Y[1333]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1334_1
  function_19 neuron1334_1 (
      .a(~input_layer[567]),
      .b(input_layer[1251]),
      .c(input_layer[780]),
      .d(input_layer[1956]),
      .y(Y[1334]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_297 for neuron1335_1
  function_297 neuron1335_1 (
      .a(input_layer[720]),
      .b(~input_layer[482]),
      .c(input_layer[1992]),
      .d(~input_layer[1078]),
      .e(~input_layer[1817]),
      .y(Y[1335]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_352 for neuron1336_1
  function_352 neuron1336_1 (
      .a(~input_layer[1504]),
      .b(input_layer[126]),
      .c(input_layer[1409]),
      .d(~input_layer[632]),
      .e(input_layer[761]),
      .f(~input_layer[603]),
      .y(Y[1336]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1337_1
  function_5 neuron1337_1 (
      .a(input_layer[681]),
      .b(~input_layer[1243]),
      .y(Y[1337]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_353 for neuron1338_1
  function_353 neuron1338_1 (
      .a(~input_layer[1694]),
      .b(input_layer[1108]),
      .c(~input_layer[693]),
      .d(~input_layer[1341]),
      .e(~input_layer[1747]),
      .f(input_layer[783]),
      .y(Y[1338]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1339_1
  function_188 neuron1339_1 (
      .a(~input_layer[746]),
      .b(input_layer[1363]),
      .c(input_layer[1438]),
      .d(input_layer[270]),
      .e(~input_layer[1780]),
      .f(input_layer[419]),
      .y(Y[1339]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1340_1
  function_26 neuron1340_1 (
      .a(~input_layer[1890]),
      .b(~input_layer[2004]),
      .y(Y[1340]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_354 for neuron1341_1
  function_354 neuron1341_1 (
      .a(~input_layer[2213]),
      .b(input_layer[296]),
      .c(input_layer[293]),
      .d(input_layer[647]),
      .e(~input_layer[2150]),
      .f(~input_layer[2196]),
      .y(Y[1341]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1342_1
  function_56 neuron1342_1 (
      .a(~input_layer[779]),
      .b(input_layer[1402]),
      .c(~input_layer[704]),
      .d(~input_layer[1005]),
      .e(input_layer[412]),
      .y(Y[1342]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_355 for neuron1343_1
  function_355 neuron1343_1 (
      .a(~input_layer[1839]),
      .b(input_layer[1543]),
      .c(~input_layer[798]),
      .d(~input_layer[454]),
      .e(~input_layer[799]),
      .f(~input_layer[1261]),
      .y(Y[1343]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1344_1
  function_120 neuron1344_1 (
      .a(input_layer[946]),
      .b(~input_layer[559]),
      .c(input_layer[231]),
      .d(input_layer[986]),
      .e(~input_layer[2008]),
      .f(~input_layer[2335]),
      .y(Y[1344]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1345_1
  function_154 neuron1345_1 (
      .a(input_layer[1317]),
      .b(input_layer[688]),
      .c(input_layer[1388]),
      .d(~input_layer[1493]),
      .e(input_layer[1327]),
      .y(Y[1345]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1346_1
  function_67 neuron1346_1 (
      .a(input_layer[1014]),
      .b(~input_layer[952]),
      .c(input_layer[1684]),
      .d(input_layer[2153]),
      .e(~input_layer[1047]),
      .y(Y[1346]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1347_1
  function_32 neuron1347_1 (
      .a(~input_layer[1128]),
      .b(input_layer[1251]),
      .c(input_layer[366]),
      .d(~input_layer[688]),
      .y(Y[1347]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1348_1
  function_95 neuron1348_1 (
      .a(~input_layer[1446]),
      .b(input_layer[1353]),
      .c(~input_layer[558]),
      .d(~input_layer[1820]),
      .y(Y[1348]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1349_1
  function_90 neuron1349_1 (
      .a(~input_layer[293]),
      .b(input_layer[1788]),
      .c(~input_layer[1105]),
      .d(~input_layer[1370]),
      .e(~input_layer[1089]),
      .y(Y[1349]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron1350_1
  function_61 neuron1350_1 (
      .a(~input_layer[981]),
      .b(input_layer[1255]),
      .c(~input_layer[2146]),
      .d(~input_layer[2320]),
      .e(input_layer[2172]),
      .y(Y[1350]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1351_1
  function_11 neuron1351_1 (
      .a(input_layer[407]),
      .b(input_layer[1698]),
      .c(input_layer[190]),
      .d(input_layer[536]),
      .y(Y[1351]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_164 for neuron1352_1
  function_164 neuron1352_1 (
      .a(~input_layer[1696]),
      .b(input_layer[1555]),
      .c(input_layer[2332]),
      .d(input_layer[1925]),
      .e(input_layer[1792]),
      .y(Y[1352]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1353_1
  function_14 neuron1353_1 (
      .a(~input_layer[635]),
      .b(~input_layer[2309]),
      .c(input_layer[1127]),
      .d(~input_layer[2088]),
      .e(~input_layer[1635]),
      .y(Y[1353]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_356 for neuron1354_1
  function_356 neuron1354_1 (
      .a(input_layer[1028]),
      .b(input_layer[875]),
      .c(~input_layer[1629]),
      .d(~input_layer[1920]),
      .e(input_layer[856]),
      .f(input_layer[536]),
      .y(Y[1354]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1355_1
  function_18 neuron1355_1 (
      .a(~input_layer[1985]),
      .b(~input_layer[1655]),
      .c(~input_layer[1775]),
      .d(~input_layer[2112]),
      .e(input_layer[390]),
      .y(Y[1355]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1356_1
  function_12 neuron1356_1 (
      .a(~input_layer[1659]),
      .b(~input_layer[1564]),
      .c(~input_layer[1727]),
      .y(Y[1356]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_357 for neuron1357_1
  function_357 neuron1357_1 (
      .a(~input_layer[1752]),
      .b(~input_layer[1886]),
      .c(input_layer[932]),
      .d(input_layer[1328]),
      .e(input_layer[2304]),
      .f(~input_layer[2151]),
      .y(Y[1357]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1358_1
  function_14 neuron1358_1 (
      .a(~input_layer[942]),
      .b(~input_layer[1595]),
      .c(~input_layer[1425]),
      .d(~input_layer[1259]),
      .e(~input_layer[343]),
      .y(Y[1358]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron1359_1
  function_192 neuron1359_1 (
      .a(~input_layer[442]),
      .b(~input_layer[2201]),
      .c(~input_layer[1410]),
      .d(~input_layer[1371]),
      .e(input_layer[771]),
      .f(~input_layer[2281]),
      .y(Y[1359]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1360_1
  function_11 neuron1360_1 (
      .a(input_layer[1239]),
      .b(input_layer[1651]),
      .c(input_layer[1955]),
      .d(~input_layer[1381]),
      .y(Y[1360]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1361_1
  function_3 neuron1361_1 (
      .a(input_layer[2238]),
      .b(input_layer[1522]),
      .c(input_layer[2142]),
      .d(~input_layer[1994]),
      .e(~input_layer[1057]),
      .y(Y[1361]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1362_1
  function_16 neuron1362_1 (
      .a(input_layer[234]),
      .b(~input_layer[1036]),
      .c(input_layer[1794]),
      .y(Y[1362]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1363_1
  function_56 neuron1363_1 (
      .a(~input_layer[1589]),
      .b(input_layer[1971]),
      .c(~input_layer[927]),
      .d(input_layer[1032]),
      .e(~input_layer[557]),
      .y(Y[1363]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1364_1
  function_44 neuron1364_1 (
      .a(input_layer[1629]),
      .b(input_layer[1499]),
      .c(~input_layer[693]),
      .y(Y[1364]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_341 for neuron1365_1
  function_341 neuron1365_1 (
      .a(input_layer[1184]),
      .b(input_layer[1679]),
      .c(~input_layer[880]),
      .d(~input_layer[560]),
      .e(~input_layer[1522]),
      .f(input_layer[577]),
      .y(Y[1365]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1366_1
  function_135 neuron1366_1 (
      .a(~input_layer[1219]),
      .b(input_layer[2070]),
      .c(~input_layer[308]),
      .d(input_layer[573]),
      .e(input_layer[1907]),
      .y(Y[1366]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_292 for neuron1367_1
  function_292 neuron1367_1 (
      .a(~input_layer[351]),
      .b(~input_layer[148]),
      .c(input_layer[1240]),
      .d(~input_layer[1172]),
      .e(input_layer[938]),
      .f(input_layer[1508]),
      .y(Y[1367]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1368_1
  function_67 neuron1368_1 (
      .a(input_layer[409]),
      .b(~input_layer[1383]),
      .c(input_layer[976]),
      .d(input_layer[352]),
      .e(~input_layer[2075]),
      .y(Y[1368]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1369_1
  function_20 neuron1369_1 (
      .a(input_layer[881]),
      .b(input_layer[874]),
      .c(input_layer[2244]),
      .d(input_layer[1327]),
      .e(input_layer[414]),
      .f(~input_layer[886]),
      .y(Y[1369]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1370_1
  function_12 neuron1370_1 (
      .a(~input_layer[1540]),
      .b(~input_layer[1080]),
      .c(~input_layer[324]),
      .y(Y[1370]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1371_1
  function_100 neuron1371_1 (
      .a(input_layer[868]),
      .b(input_layer[1291]),
      .c(~input_layer[1804]),
      .y(Y[1371]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1372_1
  function_31 neuron1372_1 (
      .a(input_layer[735]),
      .b(input_layer[1484]),
      .c(input_layer[575]),
      .d(input_layer[874]),
      .e(input_layer[2242]),
      .f(~input_layer[719]),
      .y(Y[1372]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron1373_1
  function_248 neuron1373_1 (
      .a(input_layer[523]),
      .b(~input_layer[858]),
      .c(~input_layer[215]),
      .d(~input_layer[118]),
      .e(input_layer[509]),
      .f(input_layer[1853]),
      .y(Y[1373]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1374_1
  function_107 neuron1374_1 (
      .a(input_layer[1228]),
      .b(~input_layer[2299]),
      .c(~input_layer[879]),
      .d(input_layer[712]),
      .y(Y[1374]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron1375_1
  function_133 neuron1375_1 (
      .a(~input_layer[1293]),
      .b(input_layer[1166]),
      .c(~input_layer[1771]),
      .d(input_layer[1009]),
      .e(input_layer[1073]),
      .y(Y[1375]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1376_1
  function_45 neuron1376_1 (
      .a(~input_layer[554]),
      .b(input_layer[1151]),
      .c(~input_layer[1843]),
      .d(~input_layer[2253]),
      .e(~input_layer[419]),
      .f(~input_layer[992]),
      .y(Y[1376]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_358 for neuron1377_1
  function_358 neuron1377_1 (
      .a(~input_layer[2225]),
      .b(~input_layer[2203]),
      .c(input_layer[482]),
      .d(input_layer[1575]),
      .e(input_layer[374]),
      .f(~input_layer[2057]),
      .y(Y[1377]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1378_1
  function_19 neuron1378_1 (
      .a(~input_layer[1921]),
      .b(~input_layer[2118]),
      .c(input_layer[2324]),
      .d(input_layer[1186]),
      .y(Y[1378]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_359 for neuron1379_1
  function_359 neuron1379_1 (
      .a(~input_layer[1218]),
      .b(~input_layer[1696]),
      .c(input_layer[1099]),
      .d(input_layer[1392]),
      .e(~input_layer[1604]),
      .f(~input_layer[1458]),
      .y(Y[1379]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1380_1
  function_125 neuron1380_1 (
      .a(~input_layer[463]),
      .b(~input_layer[359]),
      .c(input_layer[1306]),
      .d(input_layer[962]),
      .e(~input_layer[1674]),
      .y(Y[1380]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1381_1
  function_10 neuron1381_1 (
      .a(input_layer[2131]),
      .b(input_layer[1055]),
      .c(~input_layer[1879]),
      .d(~input_layer[379]),
      .y(Y[1381]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1382_1
  function_53 neuron1382_1 (
      .a(input_layer[1538]),
      .b(input_layer[268]),
      .c(~input_layer[953]),
      .d(input_layer[1036]),
      .e(input_layer[2027]),
      .y(Y[1382]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron1383_1
  function_192 neuron1383_1 (
      .a(~input_layer[314]),
      .b(~input_layer[226]),
      .c(~input_layer[1519]),
      .d(input_layer[712]),
      .e(input_layer[1255]),
      .f(~input_layer[1084]),
      .y(Y[1383]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1384_1
  function_25 neuron1384_1 (
      .a(input_layer[2063]),
      .b(input_layer[1189]),
      .c(input_layer[2211]),
      .d(input_layer[2045]),
      .e(input_layer[1884]),
      .y(Y[1384]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1385_1
  function_72 neuron1385_1 (
      .a(~input_layer[821]),
      .b(~input_layer[1185]),
      .c(input_layer[1799]),
      .d(~input_layer[692]),
      .e(input_layer[414]),
      .y(Y[1385]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_360 for neuron1386_1
  function_360 neuron1386_1 (
      .a(~input_layer[579]),
      .b(input_layer[930]),
      .c(~input_layer[954]),
      .d(~input_layer[1124]),
      .e(input_layer[874]),
      .f(~input_layer[1241]),
      .y(Y[1386]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1387_1
  function_67 neuron1387_1 (
      .a(input_layer[1584]),
      .b(input_layer[1522]),
      .c(input_layer[1447]),
      .d(~input_layer[1866]),
      .e(input_layer[392]),
      .y(Y[1387]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1388_1
  function_25 neuron1388_1 (
      .a(input_layer[1454]),
      .b(input_layer[1997]),
      .c(input_layer[1670]),
      .d(input_layer[1074]),
      .e(input_layer[1492]),
      .y(Y[1388]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1389_1
  function_11 neuron1389_1 (
      .a(input_layer[1187]),
      .b(input_layer[1740]),
      .c(input_layer[2310]),
      .d(input_layer[432]),
      .y(Y[1389]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1390_1
  function_100 neuron1390_1 (
      .a(input_layer[990]),
      .b(~input_layer[403]),
      .c(~input_layer[1618]),
      .y(Y[1390]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1391] = 1'b1;

  // instantiate function_92 for neuron1392_1
  function_92 neuron1392_1 (
      .a(~input_layer[2142]),
      .b(input_layer[1675]),
      .c(input_layer[1466]),
      .d(input_layer[2151]),
      .y(Y[1392]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1393_1
  function_32 neuron1393_1 (
      .a(input_layer[740]),
      .b(~input_layer[218]),
      .c(input_layer[1875]),
      .d(~input_layer[963]),
      .y(Y[1393]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1394_1
  function_40 neuron1394_1 (
      .a(~input_layer[1698]),
      .b(~input_layer[1083]),
      .c(~input_layer[1938]),
      .d(~input_layer[136]),
      .e(~input_layer[1174]),
      .f(~input_layer[1717]),
      .y(Y[1394]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_361 for neuron1395_1
  function_361 neuron1395_1 (
      .a(input_layer[1996]),
      .b(input_layer[196]),
      .c(input_layer[1742]),
      .d(~input_layer[2307]),
      .e(input_layer[1440]),
      .f(input_layer[41]),
      .y(Y[1395]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1396_1
  function_154 neuron1396_1 (
      .a(input_layer[917]),
      .b(input_layer[787]),
      .c(~input_layer[1353]),
      .d(~input_layer[545]),
      .e(input_layer[2114]),
      .y(Y[1396]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_267 for neuron1397_1
  function_267 neuron1397_1 (
      .a(input_layer[1256]),
      .b(~input_layer[887]),
      .c(input_layer[2006]),
      .d(~input_layer[2129]),
      .e(~input_layer[718]),
      .f(input_layer[1228]),
      .y(Y[1397]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_159 for neuron1398_1
  function_159 neuron1398_1 (
      .a(~input_layer[1038]),
      .b(input_layer[1694]),
      .c(input_layer[1163]),
      .d(input_layer[183]),
      .e(input_layer[1728]),
      .f(input_layer[1581]),
      .y(Y[1398]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1399_1
  function_107 neuron1399_1 (
      .a(~input_layer[1802]),
      .b(input_layer[684]),
      .c(~input_layer[1427]),
      .d(~input_layer[887]),
      .y(Y[1399]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1400_1
  function_3 neuron1400_1 (
      .a(input_layer[1714]),
      .b(input_layer[834]),
      .c(input_layer[190]),
      .d(input_layer[536]),
      .e(input_layer[526]),
      .y(Y[1400]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1401_1
  function_26 neuron1401_1 (
      .a(~input_layer[1164]),
      .b(input_layer[2044]),
      .y(Y[1401]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_212 for neuron1402_1
  function_212 neuron1402_1 (
      .a(input_layer[1607]),
      .b(~input_layer[1210]),
      .c(input_layer[583]),
      .d(input_layer[1748]),
      .e(input_layer[1931]),
      .f(~input_layer[13]),
      .y(Y[1402]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1403_1
  function_107 neuron1403_1 (
      .a(~input_layer[889]),
      .b(~input_layer[1106]),
      .c(input_layer[1137]),
      .d(input_layer[219]),
      .y(Y[1403]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1404_1
  function_14 neuron1404_1 (
      .a(~input_layer[1875]),
      .b(~input_layer[1949]),
      .c(input_layer[549]),
      .d(~input_layer[1448]),
      .e(input_layer[1195]),
      .y(Y[1404]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1405_1
  function_18 neuron1405_1 (
      .a(~input_layer[517]),
      .b(~input_layer[1661]),
      .c(input_layer[1221]),
      .d(~input_layer[699]),
      .e(input_layer[1228]),
      .y(Y[1405]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1406_1
  function_10 neuron1406_1 (
      .a(input_layer[1540]),
      .b(~input_layer[978]),
      .c(input_layer[715]),
      .d(input_layer[1640]),
      .y(Y[1406]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1407_1
  function_54 neuron1407_1 (
      .a(input_layer[948]),
      .b(input_layer[579]),
      .c(input_layer[990]),
      .d(input_layer[2313]),
      .e(input_layer[104]),
      .f(input_layer[155]),
      .y(Y[1407]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_362 for neuron1408_1
  function_362 neuron1408_1 (
      .a(~input_layer[1379]),
      .b(~input_layer[2082]),
      .c(~input_layer[119]),
      .d(input_layer[928]),
      .e(input_layer[1691]),
      .f(~input_layer[2235]),
      .y(Y[1408]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1409_1
  function_67 neuron1409_1 (
      .a(input_layer[1362]),
      .b(~input_layer[1221]),
      .c(input_layer[792]),
      .d(input_layer[1176]),
      .e(~input_layer[1659]),
      .y(Y[1409]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron1410_1
  function_202 neuron1410_1 (
      .a(~input_layer[1999]),
      .b(input_layer[2240]),
      .c(~input_layer[1284]),
      .d(input_layer[1790]),
      .e(input_layer[684]),
      .y(Y[1410]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1411_1
  function_25 neuron1411_1 (
      .a(input_layer[1650]),
      .b(input_layer[1573]),
      .c(input_layer[1443]),
      .d(~input_layer[639]),
      .e(input_layer[805]),
      .y(Y[1411]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1412_1
  function_11 neuron1412_1 (
      .a(input_layer[614]),
      .b(input_layer[871]),
      .c(input_layer[1150]),
      .d(input_layer[1115]),
      .y(Y[1412]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1413_1
  function_18 neuron1413_1 (
      .a(~input_layer[836]),
      .b(~input_layer[237]),
      .c(~input_layer[918]),
      .d(input_layer[1116]),
      .e(~input_layer[844]),
      .y(Y[1413]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_363 for neuron1414_1
  function_363 neuron1414_1 (
      .a(~input_layer[1803]),
      .b(input_layer[997]),
      .c(~input_layer[1161]),
      .d(input_layer[1012]),
      .e(~input_layer[1326]),
      .f(input_layer[2272]),
      .y(Y[1414]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1415_1
  function_64 neuron1415_1 (
      .a(input_layer[664]),
      .b(input_layer[485]),
      .c(~input_layer[974]),
      .d(input_layer[653]),
      .e(~input_layer[189]),
      .y(Y[1415]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1416_1
  function_44 neuron1416_1 (
      .a(~input_layer[1110]),
      .b(input_layer[1746]),
      .c(~input_layer[343]),
      .y(Y[1416]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_364 for neuron1417_1
  function_364 neuron1417_1 (
      .a(~input_layer[985]),
      .b(input_layer[350]),
      .c(input_layer[1435]),
      .d(~input_layer[1445]),
      .e(~input_layer[1313]),
      .f(input_layer[1170]),
      .y(Y[1417]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron1418_1
  function_115 neuron1418_1 (
      .a(input_layer[814]),
      .b(input_layer[943]),
      .c(~input_layer[1827]),
      .d(input_layer[592]),
      .e(input_layer[1434]),
      .y(Y[1418]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1419_1
  function_11 neuron1419_1 (
      .a(input_layer[1653]),
      .b(input_layer[1577]),
      .c(input_layer[743]),
      .d(input_layer[1509]),
      .y(Y[1419]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron1420_1
  function_117 neuron1420_1 (
      .a(~input_layer[2221]),
      .b(~input_layer[234]),
      .c(~input_layer[2315]),
      .d(input_layer[1498]),
      .e(input_layer[583]),
      .f(~input_layer[632]),
      .y(Y[1420]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1421_1
  function_72 neuron1421_1 (
      .a(~input_layer[709]),
      .b(~input_layer[1882]),
      .c(input_layer[1771]),
      .d(input_layer[1118]),
      .e(~input_layer[1528]),
      .y(Y[1421]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1422_1
  function_45 neuron1422_1 (
      .a(~input_layer[453]),
      .b(input_layer[1392]),
      .c(~input_layer[1910]),
      .d(~input_layer[1086]),
      .e(~input_layer[777]),
      .f(~input_layer[558]),
      .y(Y[1422]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron1423_1
  function_61 neuron1423_1 (
      .a(~input_layer[389]),
      .b(~input_layer[633]),
      .c(input_layer[2333]),
      .d(input_layer[1994]),
      .e(input_layer[508]),
      .y(Y[1423]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1424_1
  function_12 neuron1424_1 (
      .a(~input_layer[1631]),
      .b(~input_layer[1750]),
      .c(~input_layer[648]),
      .y(Y[1424]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron1425_1
  function_248 neuron1425_1 (
      .a(~input_layer[1748]),
      .b(~input_layer[1014]),
      .c(input_layer[1317]),
      .d(~input_layer[1871]),
      .e(input_layer[1982]),
      .f(~input_layer[1177]),
      .y(Y[1425]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1426_1
  function_20 neuron1426_1 (
      .a(input_layer[1798]),
      .b(input_layer[565]),
      .c(input_layer[456]),
      .d(~input_layer[784]),
      .e(input_layer[133]),
      .f(~input_layer[1026]),
      .y(Y[1426]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1427_1
  function_148 neuron1427_1 (
      .a(~input_layer[1471]),
      .b(input_layer[721]),
      .c(~input_layer[1113]),
      .d(~input_layer[1156]),
      .y(Y[1427]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1428_1
  function_113 neuron1428_1 (
      .a(input_layer[1689]),
      .b(~input_layer[531]),
      .c(input_layer[329]),
      .d(input_layer[1760]),
      .e(~input_layer[2280]),
      .f(~input_layer[596]),
      .y(Y[1428]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_332 for neuron1429_1
  function_332 neuron1429_1 (
      .a(input_layer[1585]),
      .b(input_layer[1338]),
      .c(~input_layer[2168]),
      .d(~input_layer[237]),
      .e(~input_layer[1084]),
      .f(input_layer[45]),
      .y(Y[1429]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1430_1
  function_1 neuron1430_1 (
      .a(~input_layer[1319]),
      .b(~input_layer[567]),
      .c(~input_layer[848]),
      .d(~input_layer[782]),
      .e(~input_layer[1684]),
      .f(~input_layer[2282]),
      .y(Y[1430]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_365 for neuron1431_1
  function_365 neuron1431_1 (
      .a(~input_layer[664]),
      .b(~input_layer[1131]),
      .c(input_layer[1376]),
      .d(~input_layer[739]),
      .e(input_layer[2001]),
      .y(Y[1431]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1432_1
  function_44 neuron1432_1 (
      .a(input_layer[1080]),
      .b(~input_layer[356]),
      .c(~input_layer[1673]),
      .y(Y[1432]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron1433_1
  function_253 neuron1433_1 (
      .a(~input_layer[800]),
      .b(input_layer[1870]),
      .c(input_layer[1566]),
      .d(input_layer[1367]),
      .e(input_layer[1174]),
      .y(Y[1433]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_109 for neuron1434_1
  function_109 neuron1434_1 (
      .a(input_layer[2153]),
      .b(~input_layer[1620]),
      .c(input_layer[704]),
      .d(input_layer[1341]),
      .e(input_layer[1640]),
      .f(~input_layer[1647]),
      .y(Y[1434]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1435_1
  function_113 neuron1435_1 (
      .a(input_layer[1614]),
      .b(input_layer[666]),
      .c(input_layer[800]),
      .d(~input_layer[1207]),
      .e(input_layer[1898]),
      .f(input_layer[1270]),
      .y(Y[1435]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron1436_1
  function_52 neuron1436_1 (
      .a(~input_layer[633]),
      .b(~input_layer[1563]),
      .c(input_layer[1147]),
      .d(~input_layer[1723]),
      .e(input_layer[740]),
      .y(Y[1436]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1437_1
  function_12 neuron1437_1 (
      .a(~input_layer[1163]),
      .b(input_layer[1705]),
      .c(~input_layer[1436]),
      .y(Y[1437]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1438_1
  function_148 neuron1438_1 (
      .a(~input_layer[1468]),
      .b(input_layer[1277]),
      .c(~input_layer[447]),
      .d(~input_layer[1576]),
      .y(Y[1438]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_366 for neuron1439_1
  function_366 neuron1439_1 (
      .a(~input_layer[311]),
      .b(~input_layer[1017]),
      .c(input_layer[2028]),
      .d(~input_layer[1376]),
      .e(input_layer[2325]),
      .f(input_layer[2096]),
      .y(Y[1439]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1440_1
  function_11 neuron1440_1 (
      .a(input_layer[615]),
      .b(input_layer[671]),
      .c(input_layer[416]),
      .d(input_layer[2046]),
      .y(Y[1440]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_367 for neuron1441_1
  function_367 neuron1441_1 (
      .a(~input_layer[1458]),
      .b(input_layer[413]),
      .c(input_layer[2141]),
      .d(input_layer[1401]),
      .e(~input_layer[1566]),
      .f(~input_layer[62]),
      .y(Y[1441]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1442_1
  function_76 neuron1442_1 (
      .a(~input_layer[1905]),
      .b(~input_layer[607]),
      .c(~input_layer[1095]),
      .d(~input_layer[455]),
      .e(~input_layer[924]),
      .f(input_layer[343]),
      .y(Y[1442]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1443_1
  function_10 neuron1443_1 (
      .a(input_layer[1239]),
      .b(~input_layer[533]),
      .c(input_layer[100]),
      .d(input_layer[662]),
      .y(Y[1443]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_310 for neuron1444_1
  function_310 neuron1444_1 (
      .a(~input_layer[1187]),
      .b(input_layer[1642]),
      .c(input_layer[853]),
      .d(input_layer[1985]),
      .e(input_layer[1576]),
      .f(input_layer[2250]),
      .y(Y[1444]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1445_1
  function_107 neuron1445_1 (
      .a(~input_layer[521]),
      .b(input_layer[1977]),
      .c(~input_layer[1656]),
      .d(~input_layer[1736]),
      .y(Y[1445]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_368 for neuron1446_1
  function_368 neuron1446_1 (
      .a(input_layer[1020]),
      .b(~input_layer[1040]),
      .c(input_layer[1353]),
      .d(input_layer[2261]),
      .e(~input_layer[2075]),
      .f(input_layer[2268]),
      .y(Y[1446]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_258 for neuron1447_1
  function_258 neuron1447_1 (
      .a(~input_layer[580]),
      .b(input_layer[1475]),
      .c(input_layer[1453]),
      .d(input_layer[1592]),
      .e(~input_layer[955]),
      .f(input_layer[1299]),
      .y(Y[1447]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1448_1
  function_64 neuron1448_1 (
      .a(input_layer[213]),
      .b(input_layer[398]),
      .c(~input_layer[2167]),
      .d(input_layer[437]),
      .e(~input_layer[2089]),
      .y(Y[1448]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1449_1
  function_3 neuron1449_1 (
      .a(input_layer[2154]),
      .b(input_layer[763]),
      .c(input_layer[1675]),
      .d(~input_layer[1647]),
      .e(~input_layer[1896]),
      .y(Y[1449]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_369 for neuron1450_1
  function_369 neuron1450_1 (
      .a(~input_layer[2065]),
      .b(input_layer[2115]),
      .c(~input_layer[1095]),
      .d(input_layer[2161]),
      .e(input_layer[1361]),
      .f(input_layer[594]),
      .y(Y[1450]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1451_1
  function_35 neuron1451_1 (
      .a(input_layer[1124]),
      .b(~input_layer[234]),
      .c(input_layer[953]),
      .d(~input_layer[1942]),
      .e(input_layer[2065]),
      .y(Y[1451]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1452_1
  function_26 neuron1452_1 (
      .a(~input_layer[1419]),
      .b(input_layer[1111]),
      .y(Y[1452]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1453_1
  function_146 neuron1453_1 (
      .a(input_layer[276]),
      .b(input_layer[2163]),
      .c(~input_layer[1038]),
      .d(~input_layer[1066]),
      .e(input_layer[458]),
      .y(Y[1453]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1454_1
  function_14 neuron1454_1 (
      .a(~input_layer[1990]),
      .b(~input_layer[2083]),
      .c(~input_layer[763]),
      .d(input_layer[1642]),
      .e(input_layer[193]),
      .y(Y[1454]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1455_1
  function_181 neuron1455_1 (
      .a(~input_layer[1625]),
      .b(~input_layer[2036]),
      .c(~input_layer[1510]),
      .d(~input_layer[1918]),
      .e(input_layer[2004]),
      .f(~input_layer[1814]),
      .y(Y[1455]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_170 for neuron1456_1
  function_170 neuron1456_1 (
      .a(~input_layer[1435]),
      .b(~input_layer[1542]),
      .c(~input_layer[1172]),
      .d(~input_layer[1792]),
      .e(input_layer[1112]),
      .y(Y[1456]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron1457_1
  function_34 neuron1457_1 (
      .a(input_layer[522]),
      .b(~input_layer[1538]),
      .c(input_layer[1251]),
      .d(input_layer[2327]),
      .e(input_layer[978]),
      .y(Y[1457]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_206 for neuron1458_1
  function_206 neuron1458_1 (
      .a(input_layer[1321]),
      .b(~input_layer[534]),
      .c(~input_layer[1704]),
      .d(~input_layer[1031]),
      .e(input_layer[1595]),
      .y(Y[1458]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_370 for neuron1459_1
  function_370 neuron1459_1 (
      .a(~input_layer[659]),
      .b(input_layer[2248]),
      .c(~input_layer[1534]),
      .d(input_layer[39]),
      .e(~input_layer[1839]),
      .f(input_layer[1767]),
      .y(Y[1459]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_90 for neuron1460_1
  function_90 neuron1460_1 (
      .a(~input_layer[1022]),
      .b(~input_layer[2250]),
      .c(input_layer[684]),
      .d(~input_layer[1623]),
      .e(input_layer[1563]),
      .y(Y[1460]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_371 for neuron1461_1
  function_371 neuron1461_1 (
      .a(input_layer[1665]),
      .b(input_layer[1827]),
      .c(input_layer[1473]),
      .d(~input_layer[803]),
      .e(~input_layer[593]),
      .f(input_layer[654]),
      .y(Y[1461]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1462_1
  function_298 neuron1462_1 (
      .a(input_layer[2320]),
      .b(~input_layer[1034]),
      .c(input_layer[1553]),
      .d(~input_layer[1224]),
      .e(~input_layer[1267]),
      .y(Y[1462]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1463_1
  function_107 neuron1463_1 (
      .a(~input_layer[894]),
      .b(~input_layer[913]),
      .c(input_layer[1895]),
      .d(~input_layer[671]),
      .y(Y[1463]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_257 for neuron1464_1
  function_257 neuron1464_1 (
      .a(input_layer[1628]),
      .b(~input_layer[888]),
      .c(~input_layer[856]),
      .d(~input_layer[1508]),
      .e(~input_layer[1803]),
      .y(Y[1464]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_325 for neuron1465_1
  function_325 neuron1465_1 (
      .a(input_layer[1162]),
      .b(~input_layer[971]),
      .c(input_layer[187]),
      .d(input_layer[1188]),
      .e(~input_layer[720]),
      .f(~input_layer[510]),
      .y(Y[1465]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1466_1
  function_3 neuron1466_1 (
      .a(input_layer[1782]),
      .b(input_layer[1760]),
      .c(input_layer[1436]),
      .d(input_layer[1816]),
      .e(input_layer[1965]),
      .y(Y[1466]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1467_1
  function_5 neuron1467_1 (
      .a(input_layer[1041]),
      .b(input_layer[303]),
      .y(Y[1467]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_65 for neuron1468_1
  function_65 neuron1468_1 (
      .a(~input_layer[1502]),
      .b(~input_layer[284]),
      .c(~input_layer[1626]),
      .d(input_layer[1029]),
      .e(~input_layer[822]),
      .f(~input_layer[1973]),
      .y(Y[1468]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_89 for neuron1469_1
  function_89 neuron1469_1 (
      .a(input_layer[211]),
      .b(~input_layer[2025]),
      .c(input_layer[1004]),
      .d(input_layer[134]),
      .e(~input_layer[447]),
      .f(~input_layer[291]),
      .y(Y[1469]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1470_1
  function_116 neuron1470_1 (
      .a(input_layer[2241]),
      .b(input_layer[1071]),
      .c(input_layer[327]),
      .d(~input_layer[1171]),
      .y(Y[1470]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1471_1
  function_107 neuron1471_1 (
      .a(~input_layer[1772]),
      .b(~input_layer[460]),
      .c(~input_layer[2061]),
      .d(input_layer[562]),
      .y(Y[1471]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_60 for neuron1472_1
  function_60 neuron1472_1 (
      .a(~input_layer[1573]),
      .b(input_layer[827]),
      .c(input_layer[1582]),
      .d(~input_layer[1720]),
      .e(~input_layer[1101]),
      .f(input_layer[149]),
      .y(Y[1472]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1473_1
  function_12 neuron1473_1 (
      .a(~input_layer[963]),
      .b(~input_layer[915]),
      .c(~input_layer[847]),
      .y(Y[1473]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1474_1
  function_39 neuron1474_1 (
      .a(input_layer[1858]),
      .b(input_layer[1301]),
      .c(~input_layer[1678]),
      .d(~input_layer[2000]),
      .y(Y[1474]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1475_1
  function_16 neuron1475_1 (
      .a(input_layer[484]),
      .b(input_layer[1815]),
      .c(input_layer[662]),
      .y(Y[1475]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1476_1
  function_24 neuron1476_1 (
      .a(~input_layer[1074]),
      .y(Y[1476]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_331 for neuron1477_1
  function_331 neuron1477_1 (
      .a(input_layer[599]),
      .b(input_layer[967]),
      .c(input_layer[1524]),
      .d(~input_layer[307]),
      .e(input_layer[557]),
      .y(Y[1477]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1478_1
  function_44 neuron1478_1 (
      .a(~input_layer[1231]),
      .b(~input_layer[535]),
      .c(input_layer[2173]),
      .y(Y[1478]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1479_1
  function_149 neuron1479_1 (
      .a(~input_layer[490]),
      .b(~input_layer[1950]),
      .c(~input_layer[2294]),
      .d(input_layer[1335]),
      .y(Y[1479]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_341 for neuron1480_1
  function_341 neuron1480_1 (
      .a(~input_layer[1740]),
      .b(input_layer[377]),
      .c(input_layer[1486]),
      .d(input_layer[1007]),
      .e(input_layer[1737]),
      .f(~input_layer[23]),
      .y(Y[1480]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron1481_1
  function_179 neuron1481_1 (
      .a(input_layer[1298]),
      .b(~input_layer[790]),
      .c(input_layer[152]),
      .d(~input_layer[2211]),
      .e(input_layer[1574]),
      .y(Y[1481]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_299 for neuron1482_1
  function_299 neuron1482_1 (
      .a(input_layer[2049]),
      .b(~input_layer[1908]),
      .c(input_layer[1878]),
      .d(input_layer[1018]),
      .e(input_layer[2293]),
      .f(input_layer[2175]),
      .y(Y[1482]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1483_1
  function_21 neuron1483_1 (
      .a(~input_layer[1781]),
      .b(~input_layer[1756]),
      .c(~input_layer[1501]),
      .d(input_layer[544]),
      .y(Y[1483]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_182 for neuron1484_1
  function_182 neuron1484_1 (
      .a(input_layer[912]),
      .b(~input_layer[262]),
      .c(input_layer[775]),
      .d(input_layer[476]),
      .e(~input_layer[1972]),
      .f(~input_layer[173]),
      .y(Y[1484]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron1485_1
  function_303 neuron1485_1 (
      .a(input_layer[797]),
      .b(input_layer[369]),
      .c(~input_layer[518]),
      .d(input_layer[351]),
      .e(~input_layer[791]),
      .f(input_layer[1417]),
      .y(Y[1485]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1486_1
  function_53 neuron1486_1 (
      .a(input_layer[1916]),
      .b(input_layer[2029]),
      .c(input_layer[861]),
      .d(~input_layer[1493]),
      .e(~input_layer[1952]),
      .y(Y[1486]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_79 for neuron1487_1
  function_79 neuron1487_1 (
      .a(~input_layer[1865]),
      .b(input_layer[868]),
      .c(input_layer[2173]),
      .d(input_layer[900]),
      .e(~input_layer[724]),
      .f(~input_layer[1846]),
      .y(Y[1487]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron1488_1
  function_133 neuron1488_1 (
      .a(input_layer[811]),
      .b(input_layer[1084]),
      .c(~input_layer[282]),
      .d(~input_layer[1644]),
      .e(input_layer[1782]),
      .y(Y[1488]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1489_1
  function_14 neuron1489_1 (
      .a(~input_layer[1884]),
      .b(input_layer[1291]),
      .c(~input_layer[2157]),
      .d(~input_layer[1877]),
      .e(~input_layer[587]),
      .y(Y[1489]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_174 for neuron1490_1
  function_174 neuron1490_1 (
      .a(~input_layer[2157]),
      .b(~input_layer[2090]),
      .c(input_layer[999]),
      .d(~input_layer[1921]),
      .e(input_layer[1855]),
      .f(~input_layer[132]),
      .y(Y[1490]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_197 for neuron1491_1
  function_197 neuron1491_1 (
      .a(~input_layer[433]),
      .b(~input_layer[1147]),
      .c(input_layer[105]),
      .d(input_layer[1207]),
      .e(input_layer[806]),
      .f(input_layer[1811]),
      .y(Y[1491]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron1492_1
  function_115 neuron1492_1 (
      .a(input_layer[1316]),
      .b(~input_layer[1534]),
      .c(~input_layer[866]),
      .d(input_layer[876]),
      .e(~input_layer[1950]),
      .y(Y[1492]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1493_1
  function_1 neuron1493_1 (
      .a(~input_layer[1751]),
      .b(~input_layer[766]),
      .c(~input_layer[1320]),
      .d(input_layer[1987]),
      .e(~input_layer[1759]),
      .f(~input_layer[1886]),
      .y(Y[1493]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1494_1
  function_107 neuron1494_1 (
      .a(~input_layer[830]),
      .b(~input_layer[2087]),
      .c(input_layer[882]),
      .d(input_layer[2059]),
      .y(Y[1494]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1495_1
  function_72 neuron1495_1 (
      .a(~input_layer[994]),
      .b(~input_layer[1070]),
      .c(input_layer[1435]),
      .d(input_layer[1946]),
      .e(~input_layer[2149]),
      .y(Y[1495]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1496_1
  function_307 neuron1496_1 (
      .a(input_layer[1125]),
      .b(input_layer[1974]),
      .c(~input_layer[533]),
      .d(~input_layer[565]),
      .e(~input_layer[1744]),
      .y(Y[1496]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron1497_1
  function_34 neuron1497_1 (
      .a(input_layer[602]),
      .b(~input_layer[1981]),
      .c(input_layer[301]),
      .d(input_layer[2137]),
      .e(input_layer[1154]),
      .y(Y[1497]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1498_1
  function_21 neuron1498_1 (
      .a(~input_layer[541]),
      .b(~input_layer[435]),
      .c(~input_layer[1778]),
      .d(input_layer[861]),
      .y(Y[1498]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1499_1
  function_44 neuron1499_1 (
      .a(~input_layer[1917]),
      .b(input_layer[685]),
      .c(~input_layer[1288]),
      .y(Y[1499]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_372 for neuron1500_1
  function_372 neuron1500_1 (
      .a(~input_layer[1394]),
      .b(input_layer[1064]),
      .c(input_layer[309]),
      .d(input_layer[188]),
      .e(input_layer[2253]),
      .f(~input_layer[1083]),
      .y(Y[1500]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1501_1
  function_99 neuron1501_1 (
      .a(input_layer[1528]),
      .b(input_layer[1361]),
      .c(~input_layer[2150]),
      .d(input_layer[1431]),
      .e(input_layer[101]),
      .f(~input_layer[1474]),
      .y(Y[1501]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_157 for neuron1502_1
  function_157 neuron1502_1 (
      .a(~input_layer[1944]),
      .b(input_layer[119]),
      .c(~input_layer[2114]),
      .d(input_layer[1461]),
      .e(input_layer[1628]),
      .f(input_layer[442]),
      .y(Y[1502]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1503_1
  function_26 neuron1503_1 (
      .a(~input_layer[1907]),
      .b(~input_layer[752]),
      .y(Y[1503]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1504_1
  function_95 neuron1504_1 (
      .a(input_layer[2210]),
      .b(input_layer[1074]),
      .c(~input_layer[2001]),
      .d(~input_layer[1442]),
      .y(Y[1504]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1505_1
  function_18 neuron1505_1 (
      .a(~input_layer[1971]),
      .b(~input_layer[2043]),
      .c(input_layer[1812]),
      .d(~input_layer[634]),
      .e(~input_layer[1595]),
      .y(Y[1505]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_373 for neuron1506_1
  function_373 neuron1506_1 (
      .a(input_layer[833]),
      .b(~input_layer[1280]),
      .c(input_layer[1893]),
      .d(input_layer[477]),
      .e(~input_layer[302]),
      .f(input_layer[818]),
      .y(Y[1506]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1507_1
  function_154 neuron1507_1 (
      .a(input_layer[571]),
      .b(input_layer[1502]),
      .c(~input_layer[759]),
      .d(input_layer[1904]),
      .e(~input_layer[843]),
      .y(Y[1507]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1508_1
  function_12 neuron1508_1 (
      .a(~input_layer[694]),
      .b(~input_layer[2153]),
      .c(input_layer[827]),
      .y(Y[1508]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1509_1
  function_5 neuron1509_1 (
      .a(input_layer[851]),
      .b(~input_layer[1714]),
      .y(Y[1509]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1510_1
  function_11 neuron1510_1 (
      .a(input_layer[1445]),
      .b(input_layer[1939]),
      .c(~input_layer[1140]),
      .d(input_layer[2009]),
      .y(Y[1510]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_330 for neuron1511_1
  function_330 neuron1511_1 (
      .a(input_layer[1750]),
      .b(input_layer[1365]),
      .c(input_layer[1830]),
      .d(input_layer[456]),
      .e(~input_layer[792]),
      .f(input_layer[596]),
      .y(Y[1511]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1512_1
  function_139 neuron1512_1 (
      .a(input_layer[203]),
      .b(input_layer[1816]),
      .c(input_layer[1798]),
      .d(input_layer[2126]),
      .e(input_layer[1156]),
      .y(Y[1512]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1513_1
  function_16 neuron1513_1 (
      .a(input_layer[965]),
      .b(input_layer[148]),
      .c(~input_layer[1314]),
      .y(Y[1513]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_367 for neuron1514_1
  function_367 neuron1514_1 (
      .a(input_layer[2317]),
      .b(input_layer[960]),
      .c(~input_layer[1373]),
      .d(input_layer[740]),
      .e(input_layer[113]),
      .f(~input_layer[654]),
      .y(Y[1514]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1515_1
  function_21 neuron1515_1 (
      .a(~input_layer[918]),
      .b(~input_layer[655]),
      .c(~input_layer[149]),
      .d(~input_layer[1893]),
      .y(Y[1515]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1516_1
  function_26 neuron1516_1 (
      .a(~input_layer[1065]),
      .b(~input_layer[549]),
      .y(Y[1516]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1517] = 1'b0;

  // instantiate function_16 for neuron1518_1
  function_16 neuron1518_1 (
      .a(input_layer[855]),
      .b(input_layer[112]),
      .c(~input_layer[1467]),
      .y(Y[1518]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron1519_1
  function_253 neuron1519_1 (
      .a(input_layer[384]),
      .b(~input_layer[110]),
      .c(~input_layer[2294]),
      .d(~input_layer[1763]),
      .e(input_layer[214]),
      .y(Y[1519]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1520_1
  function_1 neuron1520_1 (
      .a(~input_layer[1278]),
      .b(~input_layer[1743]),
      .c(~input_layer[687]),
      .d(input_layer[1476]),
      .e(~input_layer[2334]),
      .f(~input_layer[1973]),
      .y(Y[1520]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1521_1
  function_100 neuron1521_1 (
      .a(~input_layer[1249]),
      .b(input_layer[2244]),
      .c(input_layer[1270]),
      .y(Y[1521]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1522_1
  function_26 neuron1522_1 (
      .a(input_layer[720]),
      .b(~input_layer[1015]),
      .y(Y[1522]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1523_1
  function_231 neuron1523_1 (
      .a(~input_layer[2327]),
      .b(~input_layer[804]),
      .c(~input_layer[282]),
      .d(input_layer[445]),
      .e(~input_layer[2148]),
      .f(~input_layer[722]),
      .y(Y[1523]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1524_1
  function_125 neuron1524_1 (
      .a(~input_layer[1114]),
      .b(~input_layer[1153]),
      .c(input_layer[1735]),
      .d(input_layer[805]),
      .e(~input_layer[1294]),
      .y(Y[1524]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1525_1
  function_18 neuron1525_1 (
      .a(~input_layer[1672]),
      .b(~input_layer[1282]),
      .c(~input_layer[761]),
      .d(~input_layer[239]),
      .e(~input_layer[2254]),
      .y(Y[1525]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1526_1
  function_16 neuron1526_1 (
      .a(input_layer[1859]),
      .b(input_layer[852]),
      .c(~input_layer[1315]),
      .y(Y[1526]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1527_1
  function_12 neuron1527_1 (
      .a(~input_layer[521]),
      .b(input_layer[1974]),
      .c(~input_layer[2129]),
      .y(Y[1527]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1528_1
  function_116 neuron1528_1 (
      .a(input_layer[522]),
      .b(input_layer[1668]),
      .c(input_layer[2114]),
      .d(~input_layer[1821]),
      .y(Y[1528]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_165 for neuron1529_1
  function_165 neuron1529_1 (
      .a(~input_layer[2140]),
      .b(~input_layer[2142]),
      .c(input_layer[1191]),
      .d(~input_layer[731]),
      .e(~input_layer[1416]),
      .f(~input_layer[908]),
      .y(Y[1529]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1530_1
  function_39 neuron1530_1 (
      .a(~input_layer[1790]),
      .b(input_layer[293]),
      .c(~input_layer[2325]),
      .d(~input_layer[2177]),
      .y(Y[1530]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1531_1
  function_307 neuron1531_1 (
      .a(~input_layer[1224]),
      .b(~input_layer[107]),
      .c(input_layer[1202]),
      .d(~input_layer[1577]),
      .e(input_layer[757]),
      .y(Y[1531]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1532_1
  function_21 neuron1532_1 (
      .a(~input_layer[537]),
      .b(~input_layer[201]),
      .c(~input_layer[1574]),
      .d(input_layer[805]),
      .y(Y[1532]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_374 for neuron1533_1
  function_374 neuron1533_1 (
      .a(input_layer[998]),
      .b(input_layer[1603]),
      .c(~input_layer[1955]),
      .d(input_layer[383]),
      .e(~input_layer[2137]),
      .f(~input_layer[2043]),
      .y(Y[1533]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1534_1
  function_37 neuron1534_1 (
      .a(input_layer[1385]),
      .b(input_layer[558]),
      .c(input_layer[109]),
      .d(~input_layer[892]),
      .e(~input_layer[2143]),
      .y(Y[1534]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron1535_1
  function_133 neuron1535_1 (
      .a(input_layer[1060]),
      .b(~input_layer[1975]),
      .c(~input_layer[1667]),
      .d(input_layer[2042]),
      .e(~input_layer[486]),
      .y(Y[1535]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1536_1
  function_26 neuron1536_1 (
      .a(~input_layer[2004]),
      .b(~input_layer[738]),
      .y(Y[1536]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1537_1
  function_40 neuron1537_1 (
      .a(~input_layer[1796]),
      .b(~input_layer[1861]),
      .c(~input_layer[2114]),
      .d(~input_layer[268]),
      .e(~input_layer[103]),
      .f(input_layer[783]),
      .y(Y[1537]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1538_1
  function_107 neuron1538_1 (
      .a(~input_layer[2240]),
      .b(input_layer[1058]),
      .c(~input_layer[316]),
      .d(~input_layer[569]),
      .y(Y[1538]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron1539_1
  function_232 neuron1539_1 (
      .a(~input_layer[1498]),
      .b(input_layer[1771]),
      .c(input_layer[497]),
      .d(input_layer[1938]),
      .e(~input_layer[482]),
      .y(Y[1539]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1540_1
  function_18 neuron1540_1 (
      .a(~input_layer[216]),
      .b(~input_layer[121]),
      .c(input_layer[1275]),
      .d(~input_layer[127]),
      .e(~input_layer[1844]),
      .y(Y[1540]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1541_1
  function_64 neuron1541_1 (
      .a(input_layer[1125]),
      .b(input_layer[1069]),
      .c(input_layer[1944]),
      .d(~input_layer[1220]),
      .e(input_layer[2286]),
      .y(Y[1541]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_375 for neuron1542_1
  function_375 neuron1542_1 (
      .a(input_layer[1884]),
      .b(~input_layer[801]),
      .c(input_layer[866]),
      .d(~input_layer[391]),
      .e(~input_layer[1346]),
      .f(input_layer[2341]),
      .y(Y[1542]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron1543_1
  function_286 neuron1543_1 (
      .a(~input_layer[1137]),
      .b(~input_layer[1155]),
      .c(input_layer[1724]),
      .d(input_layer[1359]),
      .e(input_layer[1261]),
      .y(Y[1543]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1544_1
  function_26 neuron1544_1 (
      .a(~input_layer[490]),
      .b(~input_layer[2173]),
      .y(Y[1544]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1545_1
  function_125 neuron1545_1 (
      .a(~input_layer[1532]),
      .b(input_layer[1462]),
      .c(input_layer[2286]),
      .d(~input_layer[572]),
      .e(~input_layer[2092]),
      .y(Y[1545]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_376 for neuron1546_1
  function_376 neuron1546_1 (
      .a(input_layer[203]),
      .b(~input_layer[1025]),
      .c(input_layer[1073]),
      .d(~input_layer[1252]),
      .e(~input_layer[1112]),
      .f(input_layer[1262]),
      .y(Y[1546]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1547_1
  function_181 neuron1547_1 (
      .a(~input_layer[2216]),
      .b(~input_layer[1491]),
      .c(~input_layer[1269]),
      .d(input_layer[1046]),
      .e(input_layer[404]),
      .f(~input_layer[706]),
      .y(Y[1547]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1548_1
  function_149 neuron1548_1 (
      .a(~input_layer[1281]),
      .b(~input_layer[1228]),
      .c(input_layer[1550]),
      .d(~input_layer[1234]),
      .y(Y[1548]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1549_1
  function_25 neuron1549_1 (
      .a(input_layer[2138]),
      .b(input_layer[1826]),
      .c(input_layer[2082]),
      .d(input_layer[2318]),
      .e(input_layer[1146]),
      .y(Y[1549]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1550_1
  function_1 neuron1550_1 (
      .a(~input_layer[374]),
      .b(~input_layer[212]),
      .c(input_layer[1148]),
      .d(~input_layer[881]),
      .e(~input_layer[1426]),
      .f(~input_layer[1176]),
      .y(Y[1550]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1551_1
  function_25 neuron1551_1 (
      .a(input_layer[1552]),
      .b(input_layer[1495]),
      .c(input_layer[1542]),
      .d(input_layer[598]),
      .e(input_layer[106]),
      .y(Y[1551]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_163 for neuron1552_1
  function_163 neuron1552_1 (
      .a(input_layer[1221]),
      .b(input_layer[242]),
      .c(input_layer[817]),
      .d(~input_layer[1164]),
      .e(~input_layer[1322]),
      .f(~input_layer[1600]),
      .y(Y[1552]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1553_1
  function_21 neuron1553_1 (
      .a(~input_layer[1476]),
      .b(~input_layer[1605]),
      .c(~input_layer[2235]),
      .d(~input_layer[2202]),
      .y(Y[1553]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_257 for neuron1554_1
  function_257 neuron1554_1 (
      .a(input_layer[278]),
      .b(~input_layer[853]),
      .c(input_layer[1717]),
      .d(~input_layer[691]),
      .e(input_layer[372]),
      .y(Y[1554]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1555_1
  function_11 neuron1555_1 (
      .a(input_layer[549]),
      .b(input_layer[1756]),
      .c(input_layer[1752]),
      .d(~input_layer[817]),
      .y(Y[1555]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1556_1
  function_319 neuron1556_1 (
      .a(input_layer[1245]),
      .b(input_layer[2217]),
      .c(input_layer[2327]),
      .d(~input_layer[474]),
      .e(input_layer[392]),
      .f(input_layer[1008]),
      .y(Y[1556]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1557_1
  function_35 neuron1557_1 (
      .a(~input_layer[679]),
      .b(~input_layer[523]),
      .c(input_layer[2158]),
      .d(~input_layer[1818]),
      .e(~input_layer[1986]),
      .y(Y[1557]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_377 for neuron1558_1
  function_377 neuron1558_1 (
      .a(~input_layer[1510]),
      .b(input_layer[2208]),
      .c(~input_layer[1977]),
      .d(~input_layer[652]),
      .e(~input_layer[1199]),
      .f(input_layer[401]),
      .y(Y[1558]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1559_1
  function_12 neuron1559_1 (
      .a(~input_layer[456]),
      .b(~input_layer[451]),
      .c(~input_layer[1772]),
      .y(Y[1559]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_279 for neuron1560_1
  function_279 neuron1560_1 (
      .a(input_layer[1668]),
      .b(~input_layer[524]),
      .c(input_layer[390]),
      .d(~input_layer[1277]),
      .e(input_layer[350]),
      .y(Y[1560]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1561_1
  function_21 neuron1561_1 (
      .a(~input_layer[1030]),
      .b(~input_layer[1659]),
      .c(~input_layer[2305]),
      .d(~input_layer[544]),
      .y(Y[1561]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1562_1
  function_18 neuron1562_1 (
      .a(~input_layer[988]),
      .b(~input_layer[358]),
      .c(~input_layer[1839]),
      .d(~input_layer[969]),
      .e(~input_layer[151]),
      .y(Y[1562]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1563_1
  function_76 neuron1563_1 (
      .a(~input_layer[1704]),
      .b(~input_layer[2037]),
      .c(~input_layer[1864]),
      .d(input_layer[1206]),
      .e(~input_layer[1862]),
      .f(input_layer[695]),
      .y(Y[1563]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_378 for neuron1564_1
  function_378 neuron1564_1 (
      .a(~input_layer[831]),
      .b(~input_layer[995]),
      .c(input_layer[2310]),
      .d(~input_layer[1701]),
      .e(~input_layer[540]),
      .f(~input_layer[953]),
      .y(Y[1564]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1565_1
  function_11 neuron1565_1 (
      .a(input_layer[1991]),
      .b(input_layer[1017]),
      .c(input_layer[679]),
      .d(~input_layer[1386]),
      .y(Y[1565]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_262 for neuron1566_1
  function_262 neuron1566_1 (
      .a(input_layer[1479]),
      .b(input_layer[914]),
      .c(input_layer[1701]),
      .d(~input_layer[1084]),
      .e(input_layer[593]),
      .f(input_layer[1688]),
      .y(Y[1566]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1567_1
  function_104 neuron1567_1 (
      .a(~input_layer[1410]),
      .b(input_layer[1187]),
      .c(~input_layer[1436]),
      .y(Y[1567]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1568_1
  function_21 neuron1568_1 (
      .a(~input_layer[1047]),
      .b(~input_layer[1744]),
      .c(~input_layer[215]),
      .d(~input_layer[499]),
      .y(Y[1568]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1569_1
  function_3 neuron1569_1 (
      .a(input_layer[1690]),
      .b(input_layer[1591]),
      .c(input_layer[1861]),
      .d(~input_layer[205]),
      .e(~input_layer[1389]),
      .y(Y[1569]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1570_1
  function_37 neuron1570_1 (
      .a(input_layer[1082]),
      .b(input_layer[136]),
      .c(~input_layer[407]),
      .d(~input_layer[517]),
      .e(input_layer[1946]),
      .y(Y[1570]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1571_1
  function_67 neuron1571_1 (
      .a(input_layer[1665]),
      .b(input_layer[662]),
      .c(input_layer[473]),
      .d(~input_layer[366]),
      .e(~input_layer[2114]),
      .y(Y[1571]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1572_1
  function_11 neuron1572_1 (
      .a(input_layer[591]),
      .b(input_layer[125]),
      .c(~input_layer[1302]),
      .d(~input_layer[810]),
      .y(Y[1572]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1573_1
  function_5 neuron1573_1 (
      .a(input_layer[2040]),
      .b(~input_layer[1662]),
      .y(Y[1573]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron1574_1
  function_93 neuron1574_1 (
      .a(~input_layer[484]),
      .b(~input_layer[664]),
      .c(input_layer[1130]),
      .d(~input_layer[2324]),
      .e(input_layer[2134]),
      .f(~input_layer[278]),
      .y(Y[1574]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_379 for neuron1575_1
  function_379 neuron1575_1 (
      .a(input_layer[2230]),
      .b(input_layer[992]),
      .c(~input_layer[2169]),
      .d(input_layer[315]),
      .e(input_layer[2173]),
      .f(~input_layer[1509]),
      .y(Y[1575]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1576_1
  function_26 neuron1576_1 (
      .a(~input_layer[1970]),
      .b(input_layer[379]),
      .y(Y[1576]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_380 for neuron1577_1
  function_380 neuron1577_1 (
      .a(input_layer[2033]),
      .b(~input_layer[913]),
      .c(input_layer[1350]),
      .d(~input_layer[992]),
      .e(input_layer[709]),
      .f(~input_layer[1304]),
      .y(Y[1577]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_87 for neuron1578_1
  function_87 neuron1578_1 (
      .a(input_layer[969]),
      .b(input_layer[207]),
      .c(input_layer[591]),
      .d(input_layer[2088]),
      .e(~input_layer[939]),
      .f(~input_layer[1912]),
      .y(Y[1578]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_381 for neuron1579_1
  function_381 neuron1579_1 (
      .a(input_layer[1041]),
      .b(input_layer[230]),
      .c(~input_layer[1739]),
      .d(~input_layer[614]),
      .e(input_layer[316]),
      .f(~input_layer[2178]),
      .y(Y[1579]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1580_1
  function_18 neuron1580_1 (
      .a(~input_layer[1328]),
      .b(~input_layer[709]),
      .c(~input_layer[1831]),
      .d(~input_layer[398]),
      .e(~input_layer[1512]),
      .y(Y[1580]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron1581_1
  function_33 neuron1581_1 (
      .a(~input_layer[2111]),
      .b(input_layer[1137]),
      .c(~input_layer[294]),
      .d(~input_layer[295]),
      .e(input_layer[1834]),
      .y(Y[1581]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1582_1
  function_10 neuron1582_1 (
      .a(input_layer[2288]),
      .b(input_layer[1505]),
      .c(~input_layer[792]),
      .d(input_layer[1599]),
      .y(Y[1582]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1583_1
  function_31 neuron1583_1 (
      .a(input_layer[1608]),
      .b(input_layer[1752]),
      .c(input_layer[1999]),
      .d(input_layer[1922]),
      .e(~input_layer[1553]),
      .f(input_layer[2083]),
      .y(Y[1583]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_196 for neuron1584_1
  function_196 neuron1584_1 (
      .a(input_layer[743]),
      .b(input_layer[526]),
      .c(input_layer[442]),
      .d(input_layer[589]),
      .e(input_layer[1093]),
      .f(~input_layer[712]),
      .y(Y[1584]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_84 for neuron1585_1
  function_84 neuron1585_1 (
      .a(~input_layer[1471]),
      .b(~input_layer[1910]),
      .c(input_layer[1742]),
      .d(~input_layer[1023]),
      .e(~input_layer[261]),
      .f(~input_layer[1274]),
      .y(Y[1585]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1586_1
  function_21 neuron1586_1 (
      .a(~input_layer[2159]),
      .b(~input_layer[1253]),
      .c(~input_layer[825]),
      .d(input_layer[1141]),
      .y(Y[1586]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1587_1
  function_18 neuron1587_1 (
      .a(~input_layer[2166]),
      .b(input_layer[786]),
      .c(~input_layer[1755]),
      .d(~input_layer[659]),
      .e(~input_layer[1298]),
      .y(Y[1587]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_382 for neuron1588_1
  function_382 neuron1588_1 (
      .a(~input_layer[2115]),
      .b(~input_layer[2219]),
      .c(~input_layer[313]),
      .d(input_layer[1780]),
      .e(input_layer[940]),
      .f(input_layer[1339]),
      .y(Y[1588]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1589_1
  function_107 neuron1589_1 (
      .a(~input_layer[1058]),
      .b(~input_layer[2153]),
      .c(input_layer[1793]),
      .d(~input_layer[1100]),
      .y(Y[1589]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_383 for neuron1590_1
  function_383 neuron1590_1 (
      .a(input_layer[816]),
      .b(~input_layer[659]),
      .c(input_layer[2308]),
      .d(~input_layer[459]),
      .e(input_layer[2096]),
      .f(input_layer[695]),
      .y(Y[1590]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_228 for neuron1591_1
  function_228 neuron1591_1 (
      .a(~input_layer[614]),
      .b(~input_layer[1186]),
      .c(~input_layer[2096]),
      .d(input_layer[1958]),
      .e(~input_layer[521]),
      .f(~input_layer[94]),
      .y(Y[1591]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1592_1
  function_125 neuron1592_1 (
      .a(~input_layer[1024]),
      .b(~input_layer[1120]),
      .c(input_layer[1553]),
      .d(input_layer[1826]),
      .e(input_layer[444]),
      .y(Y[1592]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1593_1
  function_11 neuron1593_1 (
      .a(input_layer[522]),
      .b(~input_layer[1266]),
      .c(input_layer[768]),
      .d(input_layer[983]),
      .y(Y[1593]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1594_1
  function_16 neuron1594_1 (
      .a(input_layer[901]),
      .b(input_layer[2153]),
      .c(input_layer[897]),
      .y(Y[1594]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1595_1
  function_10 neuron1595_1 (
      .a(input_layer[1186]),
      .b(input_layer[1944]),
      .c(~input_layer[1326]),
      .d(input_layer[1879]),
      .y(Y[1595]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1596_1
  function_16 neuron1596_1 (
      .a(input_layer[1604]),
      .b(input_layer[1550]),
      .c(input_layer[934]),
      .y(Y[1596]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1597_1
  function_149 neuron1597_1 (
      .a(~input_layer[326]),
      .b(~input_layer[2287]),
      .c(input_layer[1731]),
      .d(~input_layer[2087]),
      .y(Y[1597]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1598_1
  function_19 neuron1598_1 (
      .a(~input_layer[749]),
      .b(input_layer[1030]),
      .c(~input_layer[1788]),
      .d(input_layer[1864]),
      .y(Y[1598]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1599_1
  function_307 neuron1599_1 (
      .a(~input_layer[390]),
      .b(input_layer[814]),
      .c(~input_layer[1254]),
      .d(input_layer[1349]),
      .e(input_layer[1093]),
      .y(Y[1599]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1600_1
  function_20 neuron1600_1 (
      .a(input_layer[446]),
      .b(~input_layer[795]),
      .c(input_layer[1259]),
      .d(input_layer[1547]),
      .e(input_layer[101]),
      .f(~input_layer[1005]),
      .y(Y[1600]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron1601_1
  function_210 neuron1601_1 (
      .a(~input_layer[1416]),
      .b(input_layer[129]),
      .c(input_layer[915]),
      .d(~input_layer[1874]),
      .e(~input_layer[1873]),
      .y(Y[1601]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_150 for neuron1602_1
  function_150 neuron1602_1 (
      .a(input_layer[1692]),
      .b(input_layer[801]),
      .c(input_layer[643]),
      .d(input_layer[778]),
      .e(~input_layer[152]),
      .f(~input_layer[578]),
      .y(Y[1602]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron1603_1
  function_130 neuron1603_1 (
      .a(input_layer[735]),
      .b(~input_layer[304]),
      .c(input_layer[1106]),
      .d(input_layer[386]),
      .e(input_layer[2053]),
      .f(~input_layer[1475]),
      .y(Y[1603]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron1604_1
  function_43 neuron1604_1 (
      .a(input_layer[1118]),
      .b(~input_layer[1603]),
      .c(~input_layer[463]),
      .d(~input_layer[1980]),
      .e(input_layer[1999]),
      .y(Y[1604]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1605_1
  function_11 neuron1605_1 (
      .a(input_layer[2317]),
      .b(input_layer[1941]),
      .c(input_layer[2112]),
      .d(input_layer[625]),
      .y(Y[1605]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1606_1
  function_3 neuron1606_1 (
      .a(input_layer[1699]),
      .b(input_layer[1233]),
      .c(input_layer[2247]),
      .d(~input_layer[1899]),
      .e(input_layer[812]),
      .y(Y[1606]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_38 for neuron1607_1
  function_38 neuron1607_1 (
      .a(input_layer[2244]),
      .b(~input_layer[1492]),
      .c(input_layer[1859]),
      .d(~input_layer[1417]),
      .e(input_layer[428]),
      .f(input_layer[1082]),
      .y(Y[1607]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1608_1
  function_169 neuron1608_1 (
      .a(input_layer[1921]),
      .b(input_layer[2311]),
      .c(~input_layer[793]),
      .d(input_layer[2040]),
      .e(input_layer[1493]),
      .f(input_layer[622]),
      .y(Y[1608]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1609_1
  function_113 neuron1609_1 (
      .a(input_layer[751]),
      .b(~input_layer[784]),
      .c(input_layer[908]),
      .d(input_layer[1817]),
      .e(input_layer[1965]),
      .f(~input_layer[2064]),
      .y(Y[1609]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1610_1
  function_21 neuron1610_1 (
      .a(~input_layer[2236]),
      .b(~input_layer[1586]),
      .c(input_layer[1118]),
      .d(~input_layer[1719]),
      .y(Y[1610]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1611_1
  function_16 neuron1611_1 (
      .a(input_layer[229]),
      .b(input_layer[2300]),
      .c(input_layer[1056]),
      .y(Y[1611]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1612_1
  function_107 neuron1612_1 (
      .a(~input_layer[1494]),
      .b(input_layer[914]),
      .c(~input_layer[603]),
      .d(~input_layer[800]),
      .y(Y[1612]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_91 for neuron1613_1
  function_91 neuron1613_1 (
      .a(input_layer[1657]),
      .b(input_layer[1914]),
      .c(~input_layer[793]),
      .d(input_layer[116]),
      .e(~input_layer[1414]),
      .f(~input_layer[1093]),
      .y(Y[1613]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1614_1
  function_72 neuron1614_1 (
      .a(~input_layer[209]),
      .b(~input_layer[720]),
      .c(~input_layer[1524]),
      .d(input_layer[2247]),
      .e(input_layer[1838]),
      .y(Y[1614]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1615_1
  function_21 neuron1615_1 (
      .a(~input_layer[745]),
      .b(input_layer[705]),
      .c(~input_layer[677]),
      .d(~input_layer[1601]),
      .y(Y[1615]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_211 for neuron1616_1
  function_211 neuron1616_1 (
      .a(input_layer[742]),
      .b(~input_layer[2323]),
      .c(~input_layer[1351]),
      .d(~input_layer[2286]),
      .e(~input_layer[508]),
      .y(Y[1616]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1617_1
  function_100 neuron1617_1 (
      .a(input_layer[306]),
      .b(input_layer[1436]),
      .c(~input_layer[1903]),
      .y(Y[1617]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1618_1
  function_162 neuron1618_1 (
      .a(~input_layer[284]),
      .b(~input_layer[1336]),
      .c(~input_layer[1466]),
      .d(input_layer[612]),
      .e(input_layer[1694]),
      .y(Y[1618]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1619_1
  function_12 neuron1619_1 (
      .a(~input_layer[2304]),
      .b(input_layer[819]),
      .c(input_layer[1331]),
      .y(Y[1619]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1620_1
  function_231 neuron1620_1 (
      .a(~input_layer[1785]),
      .b(~input_layer[1827]),
      .c(input_layer[573]),
      .d(~input_layer[1940]),
      .e(~input_layer[659]),
      .f(input_layer[525]),
      .y(Y[1620]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_384 for neuron1621_1
  function_384 neuron1621_1 (
      .a(input_layer[1782]),
      .b(~input_layer[2302]),
      .c(input_layer[2025]),
      .d(~input_layer[2175]),
      .e(~input_layer[979]),
      .f(input_layer[1519]),
      .y(Y[1621]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1622_1
  function_167 neuron1622_1 (
      .a(input_layer[1138]),
      .b(~input_layer[1361]),
      .c(input_layer[567]),
      .d(~input_layer[594]),
      .e(input_layer[179]),
      .y(Y[1622]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1623_1
  function_11 neuron1623_1 (
      .a(input_layer[749]),
      .b(input_layer[2299]),
      .c(input_layer[974]),
      .d(input_layer[1342]),
      .y(Y[1623]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_385 for neuron1624_1
  function_385 neuron1624_1 (
      .a(input_layer[2247]),
      .b(~input_layer[806]),
      .c(input_layer[1072]),
      .d(~input_layer[804]),
      .e(input_layer[378]),
      .f(~input_layer[644]),
      .y(Y[1624]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1625_1
  function_107 neuron1625_1 (
      .a(~input_layer[406]),
      .b(~input_layer[405]),
      .c(~input_layer[675]),
      .d(~input_layer[2323]),
      .y(Y[1625]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1626_1
  function_4 neuron1626_1 (
      .a(input_layer[2053]),
      .b(~input_layer[1376]),
      .c(~input_layer[235]),
      .d(input_layer[351]),
      .e(input_layer[587]),
      .y(Y[1626]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_234 for neuron1627_1
  function_234 neuron1627_1 (
      .a(~input_layer[1225]),
      .b(~input_layer[135]),
      .c(~input_layer[1257]),
      .d(input_layer[1112]),
      .e(~input_layer[1903]),
      .f(~input_layer[481]),
      .y(Y[1627]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_386 for neuron1628_1
  function_386 neuron1628_1 (
      .a(~input_layer[311]),
      .b(input_layer[1228]),
      .c(input_layer[2116]),
      .d(input_layer[837]),
      .e(input_layer[1097]),
      .f(~input_layer[176]),
      .y(Y[1628]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_387 for neuron1629_1
  function_387 neuron1629_1 (
      .a(input_layer[773]),
      .b(~input_layer[397]),
      .c(input_layer[1197]),
      .d(~input_layer[1049]),
      .e(~input_layer[2010]),
      .f(~input_layer[1761]),
      .y(Y[1629]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1630_1
  function_307 neuron1630_1 (
      .a(~input_layer[2231]),
      .b(~input_layer[1205]),
      .c(input_layer[1701]),
      .d(~input_layer[1597]),
      .e(~input_layer[670]),
      .y(Y[1630]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_193 for neuron1631_1
  function_193 neuron1631_1 (
      .a(input_layer[826]),
      .b(input_layer[1694]),
      .c(input_layer[730]),
      .d(~input_layer[1061]),
      .e(~input_layer[1476]),
      .f(~input_layer[1381]),
      .y(Y[1631]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_39 for neuron1632_1
  function_39 neuron1632_1 (
      .a(input_layer[1146]),
      .b(input_layer[621]),
      .c(~input_layer[1816]),
      .d(~input_layer[619]),
      .y(Y[1632]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1633_1
  function_21 neuron1633_1 (
      .a(~input_layer[703]),
      .b(~input_layer[940]),
      .c(~input_layer[1255]),
      .d(~input_layer[1603]),
      .y(Y[1633]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_110 for neuron1634_1
  function_110 neuron1634_1 (
      .a(input_layer[409]),
      .b(~input_layer[1785]),
      .c(~input_layer[2289]),
      .d(input_layer[1476]),
      .e(~input_layer[680]),
      .f(~input_layer[1613]),
      .y(Y[1634]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_388 for neuron1635_1
  function_388 neuron1635_1 (
      .a(~input_layer[2222]),
      .b(~input_layer[973]),
      .c(input_layer[1916]),
      .d(~input_layer[877]),
      .e(input_layer[567]),
      .y(Y[1635]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_181 for neuron1636_1
  function_181 neuron1636_1 (
      .a(~input_layer[554]),
      .b(~input_layer[2000]),
      .c(input_layer[890]),
      .d(~input_layer[1907]),
      .e(~input_layer[2127]),
      .f(input_layer[2123]),
      .y(Y[1636]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1637_1
  function_5 neuron1637_1 (
      .a(input_layer[500]),
      .b(input_layer[1157]),
      .y(Y[1637]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1638_1
  function_0 neuron1638_1 (
      .a(input_layer[1547]),
      .b(~input_layer[699]),
      .c(input_layer[1266]),
      .d(input_layer[534]),
      .e(input_layer[1999]),
      .y(Y[1638]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_389 for neuron1639_1
  function_389 neuron1639_1 (
      .a(~input_layer[204]),
      .b(~input_layer[113]),
      .c(input_layer[1911]),
      .d(input_layer[781]),
      .e(input_layer[1755]),
      .f(input_layer[2044]),
      .y(Y[1639]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_390 for neuron1640_1
  function_390 neuron1640_1 (
      .a(input_layer[1978]),
      .b(input_layer[1991]),
      .c(input_layer[903]),
      .d(~input_layer[522]),
      .e(~input_layer[1207]),
      .f(~input_layer[2168]),
      .y(Y[1640]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_391 for neuron1641_1
  function_391 neuron1641_1 (
      .a(input_layer[1400]),
      .b(input_layer[318]),
      .c(~input_layer[1226]),
      .d(input_layer[1090]),
      .e(input_layer[956]),
      .y(Y[1641]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_392 for neuron1642_1
  function_392 neuron1642_1 (
      .a(input_layer[990]),
      .b(~input_layer[1460]),
      .c(input_layer[2294]),
      .d(~input_layer[775]),
      .e(input_layer[1691]),
      .f(~input_layer[361]),
      .y(Y[1642]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1643_1
  function_45 neuron1643_1 (
      .a(~input_layer[209]),
      .b(~input_layer[2217]),
      .c(~input_layer[761]),
      .d(~input_layer[264]),
      .e(input_layer[1478]),
      .f(~input_layer[1920]),
      .y(Y[1643]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_133 for neuron1644_1
  function_133 neuron1644_1 (
      .a(~input_layer[1660]),
      .b(input_layer[2307]),
      .c(input_layer[2288]),
      .d(~input_layer[1951]),
      .e(input_layer[2335]),
      .y(Y[1644]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1645_1
  function_99 neuron1645_1 (
      .a(input_layer[2222]),
      .b(input_layer[2328]),
      .c(~input_layer[1113]),
      .d(input_layer[1693]),
      .e(input_layer[329]),
      .f(input_layer[2177]),
      .y(Y[1645]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_393 for neuron1646_1
  function_393 neuron1646_1 (
      .a(input_layer[2071]),
      .b(~input_layer[199]),
      .c(input_layer[838]),
      .d(input_layer[1817]),
      .e(~input_layer[2000]),
      .f(~input_layer[1852]),
      .y(Y[1646]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_394 for neuron1647_1
  function_394 neuron1647_1 (
      .a(input_layer[1544]),
      .b(~input_layer[1966]),
      .c(~input_layer[432]),
      .d(input_layer[1895]),
      .e(~input_layer[1851]),
      .f(input_layer[1261]),
      .y(Y[1647]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1648_1
  function_104 neuron1648_1 (
      .a(input_layer[446]),
      .b(~input_layer[1818]),
      .c(~input_layer[494]),
      .y(Y[1648]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1649_1
  function_63 neuron1649_1 (
      .a(input_layer[220]),
      .b(input_layer[695]),
      .c(~input_layer[1315]),
      .d(~input_layer[1020]),
      .y(Y[1649]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_62 for neuron1650_1
  function_62 neuron1650_1 (
      .a(input_layer[1641]),
      .b(~input_layer[821]),
      .c(~input_layer[2293]),
      .d(input_layer[152]),
      .y(Y[1650]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_395 for neuron1651_1
  function_395 neuron1651_1 (
      .a(input_layer[682]),
      .b(input_layer[1442]),
      .c(input_layer[1358]),
      .d(input_layer[2240]),
      .e(~input_layer[1707]),
      .f(~input_layer[1791]),
      .y(Y[1651]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1652_1
  function_31 neuron1652_1 (
      .a(input_layer[2166]),
      .b(input_layer[312]),
      .c(input_layer[1232]),
      .d(input_layer[803]),
      .e(input_layer[288]),
      .f(~input_layer[1552]),
      .y(Y[1652]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1653_1
  function_18 neuron1653_1 (
      .a(~input_layer[745]),
      .b(~input_layer[1456]),
      .c(~input_layer[1379]),
      .d(~input_layer[1296]),
      .e(~input_layer[752]),
      .y(Y[1653]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1654_1
  function_139 neuron1654_1 (
      .a(input_layer[280]),
      .b(~input_layer[2142]),
      .c(~input_layer[1230]),
      .d(~input_layer[2110]),
      .e(~input_layer[617]),
      .y(Y[1654]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1655_1
  function_53 neuron1655_1 (
      .a(input_layer[1986]),
      .b(input_layer[1621]),
      .c(input_layer[2317]),
      .d(~input_layer[297]),
      .e(input_layer[857]),
      .y(Y[1655]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1656_1
  function_167 neuron1656_1 (
      .a(~input_layer[1380]),
      .b(input_layer[1585]),
      .c(~input_layer[2070]),
      .d(~input_layer[2293]),
      .e(input_layer[1851]),
      .y(Y[1656]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1657_1
  function_1 neuron1657_1 (
      .a(~input_layer[570]),
      .b(~input_layer[538]),
      .c(~input_layer[1914]),
      .d(~input_layer[631]),
      .e(~input_layer[1442]),
      .f(input_layer[2294]),
      .y(Y[1657]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1658_1
  function_54 neuron1658_1 (
      .a(input_layer[1159]),
      .b(input_layer[2199]),
      .c(input_layer[1083]),
      .d(input_layer[1534]),
      .e(input_layer[2093]),
      .f(~input_layer[973]),
      .y(Y[1658]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1659_1
  function_100 neuron1659_1 (
      .a(input_layer[1165]),
      .b(input_layer[1284]),
      .c(~input_layer[769]),
      .y(Y[1659]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1660_1
  function_125 neuron1660_1 (
      .a(input_layer[735]),
      .b(~input_layer[364]),
      .c(~input_layer[124]),
      .d(~input_layer[1491]),
      .e(~input_layer[2021]),
      .y(Y[1660]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1661_1
  function_24 neuron1661_1 (
      .a(input_layer[1464]),
      .y(Y[1661]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1662_1
  function_12 neuron1662_1 (
      .a(~input_layer[1618]),
      .b(~input_layer[1832]),
      .c(input_layer[798]),
      .y(Y[1662]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1663_1
  function_16 neuron1663_1 (
      .a(input_layer[1189]),
      .b(input_layer[741]),
      .c(input_layer[1437]),
      .y(Y[1663]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1664_1
  function_167 neuron1664_1 (
      .a(input_layer[1204]),
      .b(~input_layer[2156]),
      .c(~input_layer[1593]),
      .d(input_layer[261]),
      .e(~input_layer[1554]),
      .y(Y[1664]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1665_1
  function_25 neuron1665_1 (
      .a(input_layer[1296]),
      .b(input_layer[291]),
      .c(input_layer[1248]),
      .d(input_layer[464]),
      .e(input_layer[1339]),
      .y(Y[1665]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_396 for neuron1666_1
  function_396 neuron1666_1 (
      .a(~input_layer[2059]),
      .b(input_layer[1336]),
      .c(input_layer[203]),
      .d(~input_layer[1972]),
      .e(~input_layer[282]),
      .f(~input_layer[802]),
      .y(Y[1666]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_397 for neuron1667_1
  function_397 neuron1667_1 (
      .a(input_layer[1285]),
      .b(~input_layer[1002]),
      .c(input_layer[942]),
      .d(~input_layer[309]),
      .e(~input_layer[2293]),
      .f(~input_layer[965]),
      .y(Y[1667]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1668_1
  function_125 neuron1668_1 (
      .a(~input_layer[730]),
      .b(~input_layer[2005]),
      .c(input_layer[136]),
      .d(input_layer[711]),
      .e(input_layer[786]),
      .y(Y[1668]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1669_1
  function_64 neuron1669_1 (
      .a(input_layer[1504]),
      .b(input_layer[1923]),
      .c(~input_layer[1812]),
      .d(~input_layer[347]),
      .e(~input_layer[148]),
      .y(Y[1669]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1670_1
  function_1 neuron1670_1 (
      .a(~input_layer[696]),
      .b(~input_layer[1622]),
      .c(~input_layer[1004]),
      .d(input_layer[1305]),
      .e(~input_layer[1213]),
      .f(~input_layer[1177]),
      .y(Y[1670]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1671_1
  function_188 neuron1671_1 (
      .a(input_layer[389]),
      .b(~input_layer[2334]),
      .c(~input_layer[1309]),
      .d(input_layer[507]),
      .e(~input_layer[250]),
      .f(input_layer[43]),
      .y(Y[1671]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1672_1
  function_148 neuron1672_1 (
      .a(input_layer[1392]),
      .b(~input_layer[1891]),
      .c(input_layer[330]),
      .d(input_layer[1197]),
      .y(Y[1672]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1673_1
  function_5 neuron1673_1 (
      .a(input_layer[2246]),
      .b(input_layer[637]),
      .y(Y[1673]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1674_1
  function_188 neuron1674_1 (
      .a(input_layer[2024]),
      .b(~input_layer[1794]),
      .c(~input_layer[702]),
      .d(~input_layer[180]),
      .e(input_layer[163]),
      .f(~input_layer[93]),
      .y(Y[1674]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1675_1
  function_44 neuron1675_1 (
      .a(~input_layer[1702]),
      .b(input_layer[1537]),
      .c(input_layer[1375]),
      .y(Y[1675]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_334 for neuron1676_1
  function_334 neuron1676_1 (
      .a(~input_layer[2132]),
      .b(input_layer[1587]),
      .c(~input_layer[1064]),
      .d(~input_layer[608]),
      .e(input_layer[1509]),
      .f(input_layer[1089]),
      .y(Y[1676]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_149 for neuron1677_1
  function_149 neuron1677_1 (
      .a(~input_layer[959]),
      .b(input_layer[768]),
      .c(~input_layer[191]),
      .d(~input_layer[138]),
      .y(Y[1677]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_308 for neuron1678_1
  function_308 neuron1678_1 (
      .a(input_layer[396]),
      .b(~input_layer[1801]),
      .c(~input_layer[676]),
      .d(input_layer[141]),
      .e(~input_layer[272]),
      .f(input_layer[1006]),
      .y(Y[1678]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_300 for neuron1679_1
  function_300 neuron1679_1 (
      .a(input_layer[1249]),
      .b(~input_layer[1387]),
      .c(~input_layer[1293]),
      .d(input_layer[545]),
      .e(input_layer[1029]),
      .y(Y[1679]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron1680_1
  function_130 neuron1680_1 (
      .a(input_layer[1323]),
      .b(~input_layer[1062]),
      .c(input_layer[1974]),
      .d(input_layer[1053]),
      .e(input_layer[1090]),
      .f(input_layer[2282]),
      .y(Y[1680]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1681_1
  function_21 neuron1681_1 (
      .a(~input_layer[383]),
      .b(~input_layer[1706]),
      .c(input_layer[1114]),
      .d(input_layer[1198]),
      .y(Y[1681]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_398 for neuron1682_1
  function_398 neuron1682_1 (
      .a(~input_layer[1131]),
      .b(~input_layer[2003]),
      .c(~input_layer[439]),
      .d(~input_layer[1577]),
      .e(~input_layer[2089]),
      .f(~input_layer[177]),
      .y(Y[1682]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_156 for neuron1683_1
  function_156 neuron1683_1 (
      .a(~input_layer[1906]),
      .b(input_layer[2032]),
      .c(~input_layer[776]),
      .d(input_layer[1951]),
      .e(~input_layer[740]),
      .y(Y[1683]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_399 for neuron1684_1
  function_399 neuron1684_1 (
      .a(input_layer[847]),
      .b(~input_layer[1956]),
      .c(input_layer[272]),
      .d(input_layer[1639]),
      .e(~input_layer[2243]),
      .f(input_layer[138]),
      .y(Y[1684]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1685_1
  function_16 neuron1685_1 (
      .a(input_layer[1028]),
      .b(input_layer[2071]),
      .c(input_layer[937]),
      .y(Y[1685]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_400 for neuron1686_1
  function_400 neuron1686_1 (
      .a(~input_layer[1308]),
      .b(input_layer[1579]),
      .c(input_layer[1743]),
      .d(~input_layer[1498]),
      .e(~input_layer[1807]),
      .f(input_layer[1128]),
      .y(Y[1686]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_146 for neuron1687_1
  function_146 neuron1687_1 (
      .a(input_layer[1754]),
      .b(input_layer[396]),
      .c(input_layer[1281]),
      .d(input_layer[364]),
      .e(input_layer[1194]),
      .y(Y[1687]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_56 for neuron1688_1
  function_56 neuron1688_1 (
      .a(~input_layer[472]),
      .b(~input_layer[1736]),
      .c(~input_layer[1605]),
      .d(~input_layer[990]),
      .e(input_layer[1483]),
      .y(Y[1688]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1689_1
  function_3 neuron1689_1 (
      .a(input_layer[1250]),
      .b(input_layer[1577]),
      .c(~input_layer[1296]),
      .d(input_layer[2030]),
      .e(input_layer[936]),
      .y(Y[1689]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_189 for neuron1690_1
  function_189 neuron1690_1 (
      .a(input_layer[2146]),
      .b(input_layer[2153]),
      .c(~input_layer[408]),
      .d(input_layer[885]),
      .e(~input_layer[507]),
      .y(Y[1690]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_401 for neuron1691_1
  function_401 neuron1691_1 (
      .a(~input_layer[812]),
      .b(input_layer[203]),
      .c(~input_layer[2093]),
      .d(input_layer[1550]),
      .e(~input_layer[1060]),
      .f(input_layer[1292]),
      .y(Y[1691]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1692_1
  function_49 neuron1692_1 (
      .a(input_layer[1251]),
      .b(input_layer[1669]),
      .c(input_layer[365]),
      .d(input_layer[381]),
      .e(input_layer[1052]),
      .f(input_layer[1356]),
      .y(Y[1692]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_114 for neuron1693_1
  function_114 neuron1693_1 (
      .a(~input_layer[1050]),
      .b(~input_layer[111]),
      .c(input_layer[2301]),
      .d(~input_layer[319]),
      .e(~input_layer[2256]),
      .f(~input_layer[1180]),
      .y(Y[1693]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1694_1
  function_24 neuron1694_1 (
      .a(input_layer[472]),
      .y(Y[1694]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_402 for neuron1695_1
  function_402 neuron1695_1 (
      .a(~input_layer[662]),
      .b(input_layer[939]),
      .c(input_layer[2322]),
      .d(input_layer[1461]),
      .e(input_layer[2150]),
      .f(~input_layer[954]),
      .y(Y[1695]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron1696_1
  function_253 neuron1696_1 (
      .a(input_layer[1025]),
      .b(input_layer[241]),
      .c(~input_layer[1992]),
      .d(~input_layer[266]),
      .e(~input_layer[922]),
      .y(Y[1696]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1697_1
  function_14 neuron1697_1 (
      .a(~input_layer[1835]),
      .b(~input_layer[1171]),
      .c(~input_layer[985]),
      .d(~input_layer[926]),
      .e(~input_layer[1862]),
      .y(Y[1697]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1698_1
  function_231 neuron1698_1 (
      .a(~input_layer[1167]),
      .b(~input_layer[1689]),
      .c(input_layer[631]),
      .d(~input_layer[1488]),
      .e(input_layer[1372]),
      .f(input_layer[712]),
      .y(Y[1698]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_155 for neuron1699_1
  function_155 neuron1699_1 (
      .a(input_layer[910]),
      .b(~input_layer[1896]),
      .c(input_layer[427]),
      .d(input_layer[2011]),
      .e(input_layer[527]),
      .y(Y[1699]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1700_1
  function_11 neuron1700_1 (
      .a(input_layer[739]),
      .b(input_layer[636]),
      .c(input_layer[2314]),
      .d(input_layer[2116]),
      .y(Y[1700]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_403 for neuron1701_1
  function_403 neuron1701_1 (
      .a(~input_layer[877]),
      .b(~input_layer[2214]),
      .c(~input_layer[763]),
      .d(input_layer[1213]),
      .e(input_layer[1421]),
      .f(input_layer[440]),
      .y(Y[1701]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1702_1
  function_11 neuron1702_1 (
      .a(input_layer[717]),
      .b(input_layer[2145]),
      .c(~input_layer[370]),
      .d(input_layer[2036]),
      .y(Y[1702]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_404 for neuron1703_1
  function_404 neuron1703_1 (
      .a(~input_layer[1953]),
      .b(~input_layer[1616]),
      .c(~input_layer[482]),
      .d(input_layer[1260]),
      .e(~input_layer[2140]),
      .f(~input_layer[557]),
      .y(Y[1703]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1704_1
  function_10 neuron1704_1 (
      .a(input_layer[1328]),
      .b(input_layer[2312]),
      .c(~input_layer[909]),
      .d(input_layer[761]),
      .y(Y[1704]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1705_1
  function_18 neuron1705_1 (
      .a(~input_layer[2218]),
      .b(~input_layer[700]),
      .c(~input_layer[1502]),
      .d(input_layer[647]),
      .e(~input_layer[1097]),
      .y(Y[1705]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1706_1
  function_5 neuron1706_1 (
      .a(input_layer[1463]),
      .b(~input_layer[979]),
      .y(Y[1706]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1707_1
  function_162 neuron1707_1 (
      .a(~input_layer[1833]),
      .b(~input_layer[1293]),
      .c(~input_layer[1757]),
      .d(~input_layer[276]),
      .e(input_layer[596]),
      .y(Y[1707]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1708_1
  function_18 neuron1708_1 (
      .a(~input_layer[1398]),
      .b(~input_layer[1521]),
      .c(~input_layer[2303]),
      .d(~input_layer[1507]),
      .e(input_layer[2056]),
      .y(Y[1708]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron1709_1
  function_145 neuron1709_1 (
      .a(input_layer[1770]),
      .b(input_layer[1195]),
      .c(~input_layer[1877]),
      .d(input_layer[2242]),
      .e(~input_layer[1418]),
      .f(input_layer[1769]),
      .y(Y[1709]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1710_1
  function_14 neuron1710_1 (
      .a(~input_layer[1695]),
      .b(~input_layer[600]),
      .c(~input_layer[1434]),
      .d(input_layer[2328]),
      .e(~input_layer[628]),
      .y(Y[1710]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1711] = 1'b0;

  // instantiate function_44 for neuron1712_1
  function_44 neuron1712_1 (
      .a(input_layer[782]),
      .b(input_layer[609]),
      .c(~input_layer[560]),
      .y(Y[1712]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_405 for neuron1713_1
  function_405 neuron1713_1 (
      .a(~input_layer[492]),
      .b(input_layer[1784]),
      .c(~input_layer[1716]),
      .d(~input_layer[591]),
      .e(~input_layer[563]),
      .f(~input_layer[1964]),
      .y(Y[1713]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_28 for neuron1714_1
  function_28 neuron1714_1 (
      .a(input_layer[658]),
      .b(~input_layer[1720]),
      .c(input_layer[1511]),
      .d(input_layer[986]),
      .e(input_layer[707]),
      .f(~input_layer[225]),
      .y(Y[1714]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1715_1
  function_16 neuron1715_1 (
      .a(input_layer[1110]),
      .b(input_layer[1610]),
      .c(~input_layer[827]),
      .y(Y[1715]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron1716_1
  function_34 neuron1716_1 (
      .a(input_layer[1101]),
      .b(~input_layer[403]),
      .c(input_layer[2301]),
      .d(input_layer[269]),
      .e(input_layer[674]),
      .y(Y[1716]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1717_1
  function_99 neuron1717_1 (
      .a(input_layer[1079]),
      .b(input_layer[208]),
      .c(input_layer[720]),
      .d(input_layer[1779]),
      .e(~input_layer[1270]),
      .f(input_layer[329]),
      .y(Y[1717]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_406 for neuron1718_1
  function_406 neuron1718_1 (
      .a(~input_layer[221]),
      .b(input_layer[1029]),
      .c(input_layer[956]),
      .d(~input_layer[1297]),
      .e(input_layer[2336]),
      .f(input_layer[2066]),
      .y(Y[1718]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_395 for neuron1719_1
  function_395 neuron1719_1 (
      .a(input_layer[140]),
      .b(input_layer[467]),
      .c(~input_layer[1229]),
      .d(input_layer[1897]),
      .e(~input_layer[1902]),
      .f(input_layer[428]),
      .y(Y[1719]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1720_1
  function_148 neuron1720_1 (
      .a(input_layer[469]),
      .b(~input_layer[716]),
      .c(~input_layer[269]),
      .d(input_layer[499]),
      .y(Y[1720]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1721_1
  function_26 neuron1721_1 (
      .a(~input_layer[663]),
      .b(input_layer[450]),
      .y(Y[1721]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_259 for neuron1722_1
  function_259 neuron1722_1 (
      .a(input_layer[547]),
      .b(input_layer[712]),
      .c(~input_layer[514]),
      .d(~input_layer[395]),
      .e(~input_layer[953]),
      .f(~input_layer[1562]),
      .y(Y[1722]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_145 for neuron1723_1
  function_145 neuron1723_1 (
      .a(input_layer[935]),
      .b(input_layer[845]),
      .c(input_layer[2127]),
      .d(input_layer[591]),
      .e(~input_layer[741]),
      .f(input_layer[1570]),
      .y(Y[1723]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1724_1
  function_12 neuron1724_1 (
      .a(~input_layer[2228]),
      .b(~input_layer[1697]),
      .c(input_layer[1985]),
      .y(Y[1724]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_348 for neuron1725_1
  function_348 neuron1725_1 (
      .a(input_layer[1023]),
      .b(~input_layer[2307]),
      .c(input_layer[1053]),
      .d(input_layer[1182]),
      .e(input_layer[398]),
      .f(~input_layer[250]),
      .y(Y[1725]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_208 for neuron1726_1
  function_208 neuron1726_1 (
      .a(~input_layer[906]),
      .b(~input_layer[701]),
      .c(~input_layer[571]),
      .d(input_layer[1266]),
      .e(input_layer[1629]),
      .f(~input_layer[1696]),
      .y(Y[1726]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_0 for neuron1727_1
  function_0 neuron1727_1 (
      .a(input_layer[1522]),
      .b(input_layer[1694]),
      .c(input_layer[2072]),
      .d(input_layer[2075]),
      .e(input_layer[669]),
      .y(Y[1727]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1728_1
  function_107 neuron1728_1 (
      .a(~input_layer[1664]),
      .b(input_layer[913]),
      .c(~input_layer[435]),
      .d(input_layer[823]),
      .y(Y[1728]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1729_1
  function_10 neuron1729_1 (
      .a(input_layer[1196]),
      .b(input_layer[1207]),
      .c(input_layer[1545]),
      .d(~input_layer[462]),
      .y(Y[1729]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1730_1
  function_21 neuron1730_1 (
      .a(~input_layer[1447]),
      .b(~input_layer[785]),
      .c(~input_layer[1248]),
      .d(~input_layer[1343]),
      .y(Y[1730]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1731_1
  function_100 neuron1731_1 (
      .a(input_layer[2129]),
      .b(~input_layer[1505]),
      .c(input_layer[1323]),
      .y(Y[1731]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1732_1
  function_49 neuron1732_1 (
      .a(input_layer[1358]),
      .b(input_layer[1606]),
      .c(input_layer[683]),
      .d(input_layer[2128]),
      .e(~input_layer[625]),
      .f(input_layer[2075]),
      .y(Y[1732]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_283 for neuron1733_1
  function_283 neuron1733_1 (
      .a(~input_layer[1032]),
      .b(~input_layer[1128]),
      .c(~input_layer[1965]),
      .d(input_layer[1295]),
      .e(~input_layer[1146]),
      .f(~input_layer[115]),
      .y(Y[1733]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_167 for neuron1734_1
  function_167 neuron1734_1 (
      .a(~input_layer[1284]),
      .b(input_layer[1103]),
      .c(~input_layer[962]),
      .d(~input_layer[601]),
      .e(input_layer[1100]),
      .y(Y[1734]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1735_1
  function_16 neuron1735_1 (
      .a(input_layer[1921]),
      .b(input_layer[1441]),
      .c(~input_layer[806]),
      .y(Y[1735]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1736_1
  function_40 neuron1736_1 (
      .a(~input_layer[469]),
      .b(~input_layer[233]),
      .c(input_layer[826]),
      .d(~input_layer[538]),
      .e(~input_layer[272]),
      .f(~input_layer[429]),
      .y(Y[1736]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_40 for neuron1737_1
  function_40 neuron1737_1 (
      .a(~input_layer[1488]),
      .b(~input_layer[286]),
      .c(~input_layer[312]),
      .d(~input_layer[1566]),
      .e(~input_layer[159]),
      .f(input_layer[253]),
      .y(Y[1737]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1738_1
  function_125 neuron1738_1 (
      .a(~input_layer[1605]),
      .b(input_layer[1036]),
      .c(~input_layer[1636]),
      .d(~input_layer[1349]),
      .e(~input_layer[1976]),
      .y(Y[1738]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1739_1
  function_100 neuron1739_1 (
      .a(~input_layer[1390]),
      .b(input_layer[1770]),
      .c(input_layer[1414]),
      .y(Y[1739]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_404 for neuron1740_1
  function_404 neuron1740_1 (
      .a(~input_layer[948]),
      .b(~input_layer[1635]),
      .c(input_layer[371]),
      .d(~input_layer[155]),
      .e(input_layer[896]),
      .f(~input_layer[1260]),
      .y(Y[1740]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1741_1
  function_11 neuron1741_1 (
      .a(input_layer[354]),
      .b(input_layer[289]),
      .c(input_layer[1839]),
      .d(input_layer[1860]),
      .y(Y[1741]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1742_1
  function_35 neuron1742_1 (
      .a(~input_layer[1543]),
      .b(~input_layer[1956]),
      .c(~input_layer[1579]),
      .d(input_layer[978]),
      .e(input_layer[1378]),
      .y(Y[1742]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1743_1
  function_12 neuron1743_1 (
      .a(~input_layer[1497]),
      .b(~input_layer[2300]),
      .c(input_layer[1142]),
      .y(Y[1743]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_407 for neuron1744_1
  function_407 neuron1744_1 (
      .a(input_layer[775]),
      .b(~input_layer[486]),
      .c(input_layer[538]),
      .d(~input_layer[2208]),
      .e(~input_layer[834]),
      .f(~input_layer[2137]),
      .y(Y[1744]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron1745_1
  function_202 neuron1745_1 (
      .a(~input_layer[955]),
      .b(~input_layer[1195]),
      .c(input_layer[1943]),
      .d(~input_layer[1240]),
      .e(~input_layer[569]),
      .y(Y[1745]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1746_1
  function_3 neuron1746_1 (
      .a(input_layer[2067]),
      .b(input_layer[139]),
      .c(input_layer[489]),
      .d(input_layer[1141]),
      .e(~input_layer[1626]),
      .y(Y[1746]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_204 for neuron1747_1
  function_204 neuron1747_1 (
      .a(~input_layer[1770]),
      .b(input_layer[2044]),
      .c(input_layer[1409]),
      .d(~input_layer[936]),
      .e(input_layer[2079]),
      .y(Y[1747]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_307 for neuron1748_1
  function_307 neuron1748_1 (
      .a(~input_layer[457]),
      .b(input_layer[373]),
      .c(~input_layer[2051]),
      .d(~input_layer[918]),
      .e(~input_layer[547]),
      .y(Y[1748]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1749_1
  function_76 neuron1749_1 (
      .a(~input_layer[1306]),
      .b(~input_layer[1391]),
      .c(~input_layer[1133]),
      .d(~input_layer[1519]),
      .e(input_layer[958]),
      .f(input_layer[1450]),
      .y(Y[1749]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1750_1
  function_21 neuron1750_1 (
      .a(~input_layer[429]),
      .b(input_layer[1913]),
      .c(~input_layer[363]),
      .d(~input_layer[1217]),
      .y(Y[1750]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1751_1
  function_18 neuron1751_1 (
      .a(~input_layer[474]),
      .b(~input_layer[776]),
      .c(input_layer[1056]),
      .d(~input_layer[1478]),
      .e(input_layer[1051]),
      .y(Y[1751]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1752_1
  function_25 neuron1752_1 (
      .a(input_layer[302]),
      .b(input_layer[288]),
      .c(input_layer[2215]),
      .d(input_layer[764]),
      .e(input_layer[931]),
      .y(Y[1752]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1753_1
  function_16 neuron1753_1 (
      .a(input_layer[406]),
      .b(input_layer[515]),
      .c(~input_layer[471]),
      .y(Y[1753]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1754_1
  function_12 neuron1754_1 (
      .a(~input_layer[1071]),
      .b(input_layer[2047]),
      .c(~input_layer[2304]),
      .y(Y[1754]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_43 for neuron1755_1
  function_43 neuron1755_1 (
      .a(input_layer[863]),
      .b(~input_layer[1528]),
      .c(~input_layer[2155]),
      .d(~input_layer[357]),
      .e(~input_layer[1963]),
      .y(Y[1755]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron1756_1
  function_115 neuron1756_1 (
      .a(input_layer[469]),
      .b(~input_layer[780]),
      .c(input_layer[358]),
      .d(input_layer[1240]),
      .e(input_layer[320]),
      .y(Y[1756]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1757_1
  function_26 neuron1757_1 (
      .a(~input_layer[870]),
      .b(~input_layer[1966]),
      .y(Y[1757]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1758_1
  function_26 neuron1758_1 (
      .a(~input_layer[642]),
      .b(~input_layer[715]),
      .y(Y[1758]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1759_1
  function_14 neuron1759_1 (
      .a(~input_layer[1382]),
      .b(~input_layer[1474]),
      .c(~input_layer[1591]),
      .d(~input_layer[608]),
      .e(input_layer[1324]),
      .y(Y[1759]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_297 for neuron1760_1
  function_297 neuron1760_1 (
      .a(input_layer[883]),
      .b(~input_layer[1484]),
      .c(~input_layer[691]),
      .d(input_layer[179]),
      .e(input_layer[1455]),
      .y(Y[1760]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1761_1
  function_44 neuron1761_1 (
      .a(input_layer[2057]),
      .b(~input_layer[225]),
      .c(input_layer[684]),
      .y(Y[1761]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_403 for neuron1762_1
  function_403 neuron1762_1 (
      .a(~input_layer[1689]),
      .b(input_layer[1965]),
      .c(~input_layer[1377]),
      .d(input_layer[984]),
      .e(~input_layer[2092]),
      .f(~input_layer[1399]),
      .y(Y[1762]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1763_1
  function_107 neuron1763_1 (
      .a(~input_layer[2080]),
      .b(input_layer[1609]),
      .c(~input_layer[281]),
      .d(~input_layer[1085]),
      .y(Y[1763]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_350 for neuron1764_1
  function_350 neuron1764_1 (
      .a(input_layer[1060]),
      .b(~input_layer[1086]),
      .c(~input_layer[546]),
      .d(~input_layer[1939]),
      .e(~input_layer[1644]),
      .y(Y[1764]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_214 for neuron1765_1
  function_214 neuron1765_1 (
      .a(~input_layer[1408]),
      .b(input_layer[1723]),
      .c(~input_layer[1939]),
      .d(~input_layer[1268]),
      .e(input_layer[706]),
      .f(input_layer[2281]),
      .y(Y[1765]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1766_1
  function_16 neuron1766_1 (
      .a(input_layer[272]),
      .b(input_layer[2158]),
      .c(~input_layer[1390]),
      .y(Y[1766]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1767] = 1'b0;

  // instantiate function_12 for neuron1768_1
  function_12 neuron1768_1 (
      .a(~input_layer[2205]),
      .b(input_layer[636]),
      .c(~input_layer[591]),
      .y(Y[1768]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_336 for neuron1769_1
  function_336 neuron1769_1 (
      .a(input_layer[846]),
      .b(~input_layer[1903]),
      .c(input_layer[314]),
      .d(input_layer[2054]),
      .e(~input_layer[1408]),
      .f(~input_layer[1329]),
      .y(Y[1769]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1770] = 1'b1;

  // instantiate function_31 for neuron1771_1
  function_31 neuron1771_1 (
      .a(input_layer[1070]),
      .b(input_layer[278]),
      .c(input_layer[834]),
      .d(input_layer[2032]),
      .e(input_layer[129]),
      .f(input_layer[1213]),
      .y(Y[1771]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_132 for neuron1772_1
  function_132 neuron1772_1 (
      .a(~input_layer[1275]),
      .b(input_layer[747]),
      .c(input_layer[1533]),
      .d(~input_layer[2218]),
      .e(~input_layer[348]),
      .y(Y[1772]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_303 for neuron1773_1
  function_303 neuron1773_1 (
      .a(input_layer[318]),
      .b(input_layer[453]),
      .c(input_layer[1749]),
      .d(input_layer[1246]),
      .e(~input_layer[2210]),
      .f(input_layer[259]),
      .y(Y[1773]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1774_1
  function_31 neuron1774_1 (
      .a(input_layer[2233]),
      .b(input_layer[281]),
      .c(input_layer[1722]),
      .d(input_layer[2302]),
      .e(input_layer[272]),
      .f(input_layer[725]),
      .y(Y[1774]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1775_1
  function_21 neuron1775_1 (
      .a(~input_layer[530]),
      .b(~input_layer[1153]),
      .c(~input_layer[526]),
      .d(~input_layer[1144]),
      .y(Y[1775]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1776_1
  function_21 neuron1776_1 (
      .a(~input_layer[1651]),
      .b(~input_layer[1697]),
      .c(~input_layer[684]),
      .d(~input_layer[663]),
      .y(Y[1776]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1777_1
  function_21 neuron1777_1 (
      .a(~input_layer[691]),
      .b(~input_layer[847]),
      .c(~input_layer[457]),
      .d(input_layer[879]),
      .y(Y[1777]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1778_1
  function_107 neuron1778_1 (
      .a(~input_layer[890]),
      .b(~input_layer[1687]),
      .c(input_layer[392]),
      .d(input_layer[1497]),
      .y(Y[1778]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1779_1
  function_49 neuron1779_1 (
      .a(input_layer[1503]),
      .b(input_layer[1335]),
      .c(input_layer[2081]),
      .d(input_layer[586]),
      .e(input_layer[2061]),
      .f(input_layer[1846]),
      .y(Y[1779]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1780_1
  function_49 neuron1780_1 (
      .a(input_layer[1108]),
      .b(input_layer[830]),
      .c(input_layer[2229]),
      .d(input_layer[2204]),
      .e(~input_layer[1667]),
      .f(input_layer[656]),
      .y(Y[1780]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1781_1
  function_107 neuron1781_1 (
      .a(~input_layer[492]),
      .b(~input_layer[847]),
      .c(input_layer[1114]),
      .d(input_layer[194]),
      .y(Y[1781]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1782_1
  function_37 neuron1782_1 (
      .a(input_layer[982]),
      .b(~input_layer[654]),
      .c(input_layer[1424]),
      .d(input_layer[2036]),
      .e(~input_layer[1798]),
      .y(Y[1782]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_380 for neuron1783_1
  function_380 neuron1783_1 (
      .a(input_layer[835]),
      .b(input_layer[500]),
      .c(~input_layer[2234]),
      .d(input_layer[483]),
      .e(~input_layer[1072]),
      .f(~input_layer[2136]),
      .y(Y[1783]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1784_1
  function_64 neuron1784_1 (
      .a(input_layer[1982]),
      .b(input_layer[581]),
      .c(input_layer[343]),
      .d(input_layer[997]),
      .e(~input_layer[1648]),
      .y(Y[1784]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_408 for neuron1785_1
  function_408 neuron1785_1 (
      .a(input_layer[1437]),
      .b(~input_layer[2117]),
      .c(~input_layer[811]),
      .d(~input_layer[1481]),
      .e(input_layer[1678]),
      .f(~input_layer[2339]),
      .y(Y[1785]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1786_1
  function_19 neuron1786_1 (
      .a(~input_layer[1876]),
      .b(input_layer[2244]),
      .c(~input_layer[1896]),
      .d(input_layer[1644]),
      .y(Y[1786]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1787_1
  function_12 neuron1787_1 (
      .a(~input_layer[2159]),
      .b(~input_layer[127]),
      .c(~input_layer[398]),
      .y(Y[1787]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_120 for neuron1788_1
  function_120 neuron1788_1 (
      .a(input_layer[991]),
      .b(~input_layer[388]),
      .c(input_layer[1986]),
      .d(~input_layer[921]),
      .e(input_layer[280]),
      .f(input_layer[313]),
      .y(Y[1788]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_92 for neuron1789_1
  function_92 neuron1789_1 (
      .a(~input_layer[320]),
      .b(input_layer[599]),
      .c(input_layer[721]),
      .d(input_layer[1269]),
      .y(Y[1789]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1790_1
  function_116 neuron1790_1 (
      .a(input_layer[1832]),
      .b(~input_layer[1145]),
      .c(input_layer[1096]),
      .d(~input_layer[1768]),
      .y(Y[1790]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_210 for neuron1791_1
  function_210 neuron1791_1 (
      .a(input_layer[1242]),
      .b(input_layer[133]),
      .c(~input_layer[1476]),
      .d(input_layer[432]),
      .e(~input_layer[1870]),
      .y(Y[1791]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_409 for neuron1792_1
  function_409 neuron1792_1 (
      .a(input_layer[475]),
      .b(input_layer[648]),
      .c(~input_layer[2317]),
      .d(~input_layer[936]),
      .e(~input_layer[1594]),
      .f(~input_layer[2159]),
      .y(Y[1792]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1793_1
  function_76 neuron1793_1 (
      .a(~input_layer[1307]),
      .b(~input_layer[584]),
      .c(~input_layer[1423]),
      .d(input_layer[1285]),
      .e(input_layer[1890]),
      .f(~input_layer[535]),
      .y(Y[1793]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1794_1
  function_1 neuron1794_1 (
      .a(~input_layer[663]),
      .b(~input_layer[702]),
      .c(~input_layer[767]),
      .d(input_layer[1721]),
      .e(input_layer[2101]),
      .f(input_layer[24]),
      .y(Y[1794]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_144 for neuron1795_1
  function_144 neuron1795_1 (
      .a(~input_layer[1301]),
      .b(input_layer[1703]),
      .c(~input_layer[321]),
      .d(input_layer[1872]),
      .e(~input_layer[239]),
      .f(input_layer[1823]),
      .y(Y[1795]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron1796_1
  function_179 neuron1796_1 (
      .a(input_layer[2309]),
      .b(~input_layer[1705]),
      .c(input_layer[1091]),
      .d(~input_layer[137]),
      .e(input_layer[2281]),
      .y(Y[1796]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_410 for neuron1797_1
  function_410 neuron1797_1 (
      .a(~input_layer[309]),
      .b(~input_layer[227]),
      .c(input_layer[1606]),
      .d(input_layer[631]),
      .e(~input_layer[102]),
      .f(~input_layer[1327]),
      .y(Y[1797]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1798_1
  function_76 neuron1798_1 (
      .a(~input_layer[2153]),
      .b(~input_layer[683]),
      .c(~input_layer[266]),
      .d(~input_layer[1812]),
      .e(~input_layer[114]),
      .f(~input_layer[248]),
      .y(Y[1798]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_286 for neuron1799_1
  function_286 neuron1799_1 (
      .a(~input_layer[1624]),
      .b(input_layer[200]),
      .c(input_layer[2230]),
      .d(~input_layer[820]),
      .e(~input_layer[521]),
      .y(Y[1799]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1800_1
  function_11 neuron1800_1 (
      .a(input_layer[1040]),
      .b(input_layer[1032]),
      .c(input_layer[993]),
      .d(input_layer[833]),
      .y(Y[1800]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_372 for neuron1801_1
  function_372 neuron1801_1 (
      .a(~input_layer[291]),
      .b(input_layer[891]),
      .c(input_layer[985]),
      .d(input_layer[2165]),
      .e(input_layer[2330]),
      .f(~input_layer[1399]),
      .y(Y[1801]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_388 for neuron1802_1
  function_388 neuron1802_1 (
      .a(~input_layer[416]),
      .b(~input_layer[207]),
      .c(~input_layer[1051]),
      .d(input_layer[1276]),
      .e(input_layer[360]),
      .y(Y[1802]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1803_1
  function_11 neuron1803_1 (
      .a(input_layer[2209]),
      .b(input_layer[845]),
      .c(input_layer[2205]),
      .d(input_layer[1288]),
      .y(Y[1803]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_411 for neuron1804_1
  function_411 neuron1804_1 (
      .a(~input_layer[1392]),
      .b(input_layer[797]),
      .c(input_layer[801]),
      .d(~input_layer[1395]),
      .e(input_layer[731]),
      .f(~input_layer[1260]),
      .y(Y[1804]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1805_1
  function_10 neuron1805_1 (
      .a(input_layer[1906]),
      .b(input_layer[1415]),
      .c(input_layer[1538]),
      .d(~input_layer[2292]),
      .y(Y[1805]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_50 for neuron1806_1
  function_50 neuron1806_1 (
      .a(~input_layer[128]),
      .b(input_layer[616]),
      .c(~input_layer[1487]),
      .d(~input_layer[263]),
      .e(~input_layer[838]),
      .y(Y[1806]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1807_1
  function_100 neuron1807_1 (
      .a(input_layer[1156]),
      .b(~input_layer[1469]),
      .c(~input_layer[2323]),
      .y(Y[1807]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_119 for neuron1808_1
  function_119 neuron1808_1 (
      .a(input_layer[1079]),
      .b(input_layer[732]),
      .c(~input_layer[1471]),
      .d(input_layer[972]),
      .e(~input_layer[1639]),
      .f(input_layer[2000]),
      .y(Y[1808]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1809_1
  function_21 neuron1809_1 (
      .a(~input_layer[218]),
      .b(~input_layer[2207]),
      .c(input_layer[1222]),
      .d(~input_layer[675]),
      .y(Y[1809]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_175 for neuron1810_1
  function_175 neuron1810_1 (
      .a(~input_layer[1977]),
      .b(input_layer[815]),
      .c(~input_layer[1787]),
      .d(~input_layer[433]),
      .e(~input_layer[575]),
      .y(Y[1810]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_34 for neuron1811_1
  function_34 neuron1811_1 (
      .a(input_layer[1698]),
      .b(~input_layer[2130]),
      .c(input_layer[839]),
      .d(input_layer[132]),
      .e(input_layer[240]),
      .y(Y[1811]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1812_1
  function_11 neuron1812_1 (
      .a(input_layer[651]),
      .b(input_layer[1737]),
      .c(input_layer[145]),
      .d(input_layer[1771]),
      .y(Y[1812]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1813_1
  function_113 neuron1813_1 (
      .a(input_layer[2059]),
      .b(input_layer[734]),
      .c(input_layer[1521]),
      .d(~input_layer[1245]),
      .e(input_layer[1514]),
      .f(input_layer[794]),
      .y(Y[1813]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1814_1
  function_10 neuron1814_1 (
      .a(input_layer[210]),
      .b(input_layer[1386]),
      .c(~input_layer[2206]),
      .d(input_layer[1867]),
      .y(Y[1814]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_412 for neuron1815_1
  function_412 neuron1815_1 (
      .a(~input_layer[2086]),
      .b(~input_layer[1757]),
      .c(input_layer[930]),
      .d(input_layer[2303]),
      .e(~input_layer[2226]),
      .f(input_layer[2024]),
      .y(Y[1815]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1816_1
  function_16 neuron1816_1 (
      .a(input_layer[1819]),
      .b(input_layer[488]),
      .c(~input_layer[615]),
      .y(Y[1816]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1817_1
  function_107 neuron1817_1 (
      .a(~input_layer[213]),
      .b(~input_layer[1162]),
      .c(input_layer[1136]),
      .d(~input_layer[547]),
      .y(Y[1817]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1818_1
  function_26 neuron1818_1 (
      .a(~input_layer[1157]),
      .b(input_layer[823]),
      .y(Y[1818]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1819_1
  function_125 neuron1819_1 (
      .a(~input_layer[2121]),
      .b(~input_layer[441]),
      .c(input_layer[732]),
      .d(input_layer[2046]),
      .e(input_layer[1193]),
      .y(Y[1819]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1820_1
  function_139 neuron1820_1 (
      .a(input_layer[2309]),
      .b(~input_layer[810]),
      .c(input_layer[1800]),
      .d(~input_layer[941]),
      .e(~input_layer[1980]),
      .y(Y[1820]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_14 for neuron1821_1
  function_14 neuron1821_1 (
      .a(~input_layer[1228]),
      .b(~input_layer[934]),
      .c(~input_layer[440]),
      .d(~input_layer[466]),
      .e(input_layer[499]),
      .y(Y[1821]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_52 for neuron1822_1
  function_52 neuron1822_1 (
      .a(~input_layer[1035]),
      .b(input_layer[2142]),
      .c(input_layer[451]),
      .d(input_layer[435]),
      .e(input_layer[1504]),
      .y(Y[1822]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_232 for neuron1823_1
  function_232 neuron1823_1 (
      .a(input_layer[2067]),
      .b(~input_layer[1379]),
      .c(input_layer[644]),
      .d(~input_layer[1707]),
      .e(input_layer[1348]),
      .y(Y[1823]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_53 for neuron1824_1
  function_53 neuron1824_1 (
      .a(input_layer[1233]),
      .b(~input_layer[2078]),
      .c(input_layer[1690]),
      .d(input_layer[1747]),
      .e(input_layer[641]),
      .y(Y[1824]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_413 for neuron1825_1
  function_413 neuron1825_1 (
      .a(~input_layer[1054]),
      .b(~input_layer[2112]),
      .c(input_layer[1999]),
      .d(~input_layer[428]),
      .e(input_layer[2137]),
      .f(input_layer[1848]),
      .y(Y[1825]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_414 for neuron1826_1
  function_414 neuron1826_1 (
      .a(~input_layer[2219]),
      .b(~input_layer[1113]),
      .c(input_layer[1658]),
      .d(~input_layer[1227]),
      .e(input_layer[298]),
      .f(~input_layer[1074]),
      .y(Y[1826]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1827_1
  function_11 neuron1827_1 (
      .a(input_layer[386]),
      .b(input_layer[680]),
      .c(input_layer[1970]),
      .d(input_layer[2054]),
      .y(Y[1827]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_276 for neuron1828_1
  function_276 neuron1828_1 (
      .a(input_layer[1026]),
      .b(~input_layer[1854]),
      .c(~input_layer[1658]),
      .d(~input_layer[472]),
      .e(input_layer[908]),
      .y(Y[1828]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_135 for neuron1829_1
  function_135 neuron1829_1 (
      .a(input_layer[1468]),
      .b(~input_layer[664]),
      .c(input_layer[1667]),
      .d(input_layer[1148]),
      .e(input_layer[930]),
      .y(Y[1829]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1830_1
  function_188 neuron1830_1 (
      .a(~input_layer[615]),
      .b(input_layer[1190]),
      .c(~input_layer[602]),
      .d(~input_layer[924]),
      .e(input_layer[985]),
      .f(~input_layer[236]),
      .y(Y[1830]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_72 for neuron1831_1
  function_72 neuron1831_1 (
      .a(~input_layer[376]),
      .b(~input_layer[1741]),
      .c(~input_layer[180]),
      .d(input_layer[652]),
      .e(input_layer[768]),
      .y(Y[1831]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_415 for neuron1832_1
  function_415 neuron1832_1 (
      .a(~input_layer[1113]),
      .b(input_layer[1423]),
      .c(~input_layer[2289]),
      .d(input_layer[314]),
      .e(input_layer[1798]),
      .f(~input_layer[428]),
      .y(Y[1832]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1833_1
  function_1 neuron1833_1 (
      .a(~input_layer[697]),
      .b(~input_layer[1507]),
      .c(~input_layer[455]),
      .d(input_layer[1053]),
      .e(~input_layer[978]),
      .f(~input_layer[1784]),
      .y(Y[1833]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1834_1
  function_21 neuron1834_1 (
      .a(~input_layer[691]),
      .b(~input_layer[751]),
      .c(~input_layer[194]),
      .d(~input_layer[1517]),
      .y(Y[1834]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_262 for neuron1835_1
  function_262 neuron1835_1 (
      .a(~input_layer[1050]),
      .b(input_layer[947]),
      .c(input_layer[1950]),
      .d(input_layer[1342]),
      .e(input_layer[2012]),
      .f(~input_layer[102]),
      .y(Y[1835]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_416 for neuron1836_1
  function_416 neuron1836_1 (
      .a(~input_layer[212]),
      .b(input_layer[626]),
      .c(~input_layer[2146]),
      .d(~input_layer[1570]),
      .e(input_layer[2064]),
      .f(input_layer[1090]),
      .y(Y[1836]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_98 for neuron1837_1
  function_98 neuron1837_1 (
      .a(~input_layer[1383]),
      .b(input_layer[1032]),
      .c(~input_layer[2208]),
      .d(input_layer[1321]),
      .e(input_layer[904]),
      .y(Y[1837]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_215 for neuron1838_1
  function_215 neuron1838_1 (
      .a(input_layer[2027]),
      .b(input_layer[1474]),
      .c(input_layer[1496]),
      .d(~input_layer[1701]),
      .e(input_layer[1739]),
      .f(~input_layer[544]),
      .y(Y[1838]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_319 for neuron1839_1
  function_319 neuron1839_1 (
      .a(input_layer[2327]),
      .b(~input_layer[1118]),
      .c(input_layer[2146]),
      .d(input_layer[754]),
      .e(input_layer[1536]),
      .f(input_layer[152]),
      .y(Y[1839]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1840_1
  function_12 neuron1840_1 (
      .a(~input_layer[781]),
      .b(~input_layer[367]),
      .c(~input_layer[978]),
      .y(Y[1840]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1841_1
  function_12 neuron1841_1 (
      .a(~input_layer[1692]),
      .b(input_layer[1971]),
      .c(~input_layer[1239]),
      .y(Y[1841]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1842_1
  function_32 neuron1842_1 (
      .a(input_layer[656]),
      .b(~input_layer[889]),
      .c(~input_layer[816]),
      .d(~input_layer[1350]),
      .y(Y[1842]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1843_1
  function_67 neuron1843_1 (
      .a(input_layer[363]),
      .b(input_layer[275]),
      .c(input_layer[132]),
      .d(input_layer[1188]),
      .e(input_layer[2076]),
      .y(Y[1843]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_248 for neuron1844_1
  function_248 neuron1844_1 (
      .a(~input_layer[1378]),
      .b(~input_layer[378]),
      .c(~input_layer[226]),
      .d(~input_layer[1041]),
      .e(input_layer[1106]),
      .f(~input_layer[1389]),
      .y(Y[1844]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_417 for neuron1845_1
  function_417 neuron1845_1 (
      .a(~input_layer[872]),
      .b(input_layer[2022]),
      .c(input_layer[2296]),
      .d(~input_layer[870]),
      .e(input_layer[1886]),
      .f(input_layer[2301]),
      .y(Y[1845]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1846_1
  function_231 neuron1846_1 (
      .a(~input_layer[291]),
      .b(~input_layer[1256]),
      .c(input_layer[1975]),
      .d(~input_layer[1115]),
      .e(~input_layer[1678]),
      .f(input_layer[1167]),
      .y(Y[1846]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1847_1
  function_67 neuron1847_1 (
      .a(input_layer[1421]),
      .b(input_layer[1244]),
      .c(~input_layer[963]),
      .d(input_layer[1153]),
      .e(input_layer[376]),
      .y(Y[1847]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1848_1
  function_12 neuron1848_1 (
      .a(~input_layer[883]),
      .b(~input_layer[1961]),
      .c(~input_layer[144]),
      .y(Y[1848]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1849_1
  function_5 neuron1849_1 (
      .a(input_layer[1776]),
      .b(~input_layer[1891]),
      .y(Y[1849]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_418 for neuron1850_1
  function_418 neuron1850_1 (
      .a(~input_layer[734]),
      .b(~input_layer[362]),
      .c(~input_layer[972]),
      .d(input_layer[1710]),
      .e(input_layer[499]),
      .f(input_layer[1194]),
      .y(Y[1850]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1851_1
  function_25 neuron1851_1 (
      .a(input_layer[1948]),
      .b(input_layer[933]),
      .c(input_layer[1518]),
      .d(~input_layer[896]),
      .e(~input_layer[1806]),
      .y(Y[1851]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1852_1
  function_35 neuron1852_1 (
      .a(~input_layer[1043]),
      .b(~input_layer[1080]),
      .c(~input_layer[1046]),
      .d(~input_layer[332]),
      .e(input_layer[2193]),
      .y(Y[1852]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_201 for neuron1853_1
  function_201 neuron1853_1 (
      .a(~input_layer[1788]),
      .b(~input_layer[832]),
      .c(input_layer[2293]),
      .d(input_layer[1358]),
      .e(input_layer[1928]),
      .y(Y[1853]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1854_1
  function_5 neuron1854_1 (
      .a(input_layer[583]),
      .b(input_layer[103]),
      .y(Y[1854]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1855_1
  function_16 neuron1855_1 (
      .a(input_layer[1087]),
      .b(~input_layer[711]),
      .c(input_layer[1501]),
      .y(Y[1855]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1856_1
  function_169 neuron1856_1 (
      .a(input_layer[1770]),
      .b(input_layer[513]),
      .c(~input_layer[1884]),
      .d(~input_layer[1833]),
      .e(input_layer[1061]),
      .f(input_layer[566]),
      .y(Y[1856]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_31 for neuron1857_1
  function_31 neuron1857_1 (
      .a(input_layer[889]),
      .b(input_layer[442]),
      .c(input_layer[2248]),
      .d(input_layer[1266]),
      .e(input_layer[1668]),
      .f(input_layer[359]),
      .y(Y[1857]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1858_1
  function_21 neuron1858_1 (
      .a(~input_layer[1751]),
      .b(~input_layer[365]),
      .c(~input_layer[1399]),
      .d(~input_layer[1412]),
      .y(Y[1858]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1859_1
  function_107 neuron1859_1 (
      .a(~input_layer[1913]),
      .b(~input_layer[197]),
      .c(input_layer[615]),
      .d(input_layer[1028]),
      .y(Y[1859]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1860_1
  function_12 neuron1860_1 (
      .a(~input_layer[360]),
      .b(~input_layer[2216]),
      .c(~input_layer[1472]),
      .y(Y[1860]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1861_1
  function_67 neuron1861_1 (
      .a(input_layer[2238]),
      .b(input_layer[1169]),
      .c(~input_layer[1481]),
      .d(input_layer[2286]),
      .e(~input_layer[1484]),
      .y(Y[1861]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_253 for neuron1862_1
  function_253 neuron1862_1 (
      .a(~input_layer[1541]),
      .b(~input_layer[1185]),
      .c(input_layer[1353]),
      .d(input_layer[1563]),
      .e(~input_layer[776]),
      .y(Y[1862]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_26 for neuron1863_1
  function_26 neuron1863_1 (
      .a(~input_layer[644]),
      .b(~input_layer[1002]),
      .y(Y[1863]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1864_1
  function_25 neuron1864_1 (
      .a(input_layer[2157]),
      .b(input_layer[517]),
      .c(input_layer[143]),
      .d(~input_layer[948]),
      .e(input_layer[1601]),
      .y(Y[1864]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_410 for neuron1865_1
  function_410 neuron1865_1 (
      .a(input_layer[918]),
      .b(~input_layer[604]),
      .c(~input_layer[901]),
      .d(~input_layer[1438]),
      .e(~input_layer[611]),
      .f(~input_layer[1683]),
      .y(Y[1865]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_152 for neuron1866_1
  function_152 neuron1866_1 (
      .a(~input_layer[2052]),
      .b(input_layer[1409]),
      .c(~input_layer[920]),
      .d(input_layer[186]),
      .e(input_layer[2298]),
      .f(input_layer[320]),
      .y(Y[1866]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1867_1
  function_3 neuron1867_1 (
      .a(input_layer[685]),
      .b(input_layer[412]),
      .c(input_layer[1434]),
      .d(~input_layer[886]),
      .e(~input_layer[560]),
      .y(Y[1867]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1868_1
  function_12 neuron1868_1 (
      .a(~input_layer[107]),
      .b(~input_layer[1810]),
      .c(input_layer[1473]),
      .y(Y[1868]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1869_1
  function_35 neuron1869_1 (
      .a(~input_layer[555]),
      .b(~input_layer[1659]),
      .c(~input_layer[593]),
      .d(~input_layer[366]),
      .e(~input_layer[2016]),
      .y(Y[1869]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1870_1
  function_16 neuron1870_1 (
      .a(input_layer[898]),
      .b(input_layer[292]),
      .c(input_layer[1457]),
      .y(Y[1870]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1871_1
  function_18 neuron1871_1 (
      .a(~input_layer[1336]),
      .b(~input_layer[184]),
      .c(~input_layer[842]),
      .d(~input_layer[1921]),
      .e(~input_layer[1761]),
      .y(Y[1871]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_419 for neuron1872_1
  function_419 neuron1872_1 (
      .a(~input_layer[447]),
      .b(input_layer[1118]),
      .c(~input_layer[1086]),
      .d(~input_layer[558]),
      .e(~input_layer[1370]),
      .f(~input_layer[1679]),
      .y(Y[1872]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_24 for neuron1873_1
  function_24 neuron1873_1 (
      .a(~input_layer[1673]),
      .y(Y[1873]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_4 for neuron1874_1
  function_4 neuron1874_1 (
      .a(input_layer[1993]),
      .b(input_layer[1897]),
      .c(~input_layer[192]),
      .d(input_layer[1440]),
      .e(~input_layer[605]),
      .y(Y[1874]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_420 for neuron1875_1
  function_420 neuron1875_1 (
      .a(~input_layer[2252]),
      .b(~input_layer[971]),
      .c(input_layer[1195]),
      .d(input_layer[1583]),
      .e(input_layer[181]),
      .f(input_layer[1318]),
      .y(Y[1875]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_124 for neuron1876_1
  function_124 neuron1876_1 (
      .a(~input_layer[1357]),
      .b(input_layer[530]),
      .c(~input_layer[1854]),
      .d(input_layer[863]),
      .e(input_layer[701]),
      .f(input_layer[1873]),
      .y(Y[1876]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1877_1
  function_100 neuron1877_1 (
      .a(input_layer[1506]),
      .b(~input_layer[1296]),
      .c(~input_layer[967]),
      .y(Y[1877]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1878] = 1'b0;

  // instantiate function_146 for neuron1879_1
  function_146 neuron1879_1 (
      .a(input_layer[2239]),
      .b(~input_layer[1867]),
      .c(~input_layer[1196]),
      .d(~input_layer[1107]),
      .e(input_layer[2067]),
      .y(Y[1879]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_44 for neuron1880_1
  function_44 neuron1880_1 (
      .a(~input_layer[931]),
      .b(input_layer[877]),
      .c(input_layer[1818]),
      .y(Y[1880]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_363 for neuron1881_1
  function_363 neuron1881_1 (
      .a(input_layer[1219]),
      .b(input_layer[835]),
      .c(~input_layer[2064]),
      .d(~input_layer[2189]),
      .e(input_layer[11]),
      .f(~input_layer[72]),
      .y(Y[1881]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_76 for neuron1882_1
  function_76 neuron1882_1 (
      .a(~input_layer[1142]),
      .b(~input_layer[2212]),
      .c(~input_layer[1019]),
      .d(~input_layer[760]),
      .e(input_layer[1879]),
      .f(~input_layer[1777]),
      .y(Y[1882]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1883_1
  function_11 neuron1883_1 (
      .a(input_layer[880]),
      .b(input_layer[1584]),
      .c(~input_layer[2039]),
      .d(input_layer[2120]),
      .y(Y[1883]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1884_1
  function_107 neuron1884_1 (
      .a(~input_layer[1249]),
      .b(~input_layer[189]),
      .c(input_layer[532]),
      .d(input_layer[1804]),
      .y(Y[1884]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1885_1
  function_113 neuron1885_1 (
      .a(input_layer[1634]),
      .b(input_layer[942]),
      .c(input_layer[1673]),
      .d(input_layer[1333]),
      .e(input_layer[824]),
      .f(input_layer[1564]),
      .y(Y[1885]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1886_1
  function_162 neuron1886_1 (
      .a(~input_layer[481]),
      .b(~input_layer[1925]),
      .c(input_layer[1994]),
      .d(~input_layer[1320]),
      .e(input_layer[1392]),
      .y(Y[1886]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1887_1
  function_12 neuron1887_1 (
      .a(~input_layer[570]),
      .b(~input_layer[1704]),
      .c(input_layer[627]),
      .y(Y[1887]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_126 for neuron1888_1
  function_126 neuron1888_1 (
      .a(~input_layer[1415]),
      .b(input_layer[525]),
      .c(~input_layer[1647]),
      .d(input_layer[1612]),
      .e(input_layer[180]),
      .y(Y[1888]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1889_1
  function_18 neuron1889_1 (
      .a(~input_layer[786]),
      .b(~input_layer[693]),
      .c(~input_layer[1668]),
      .d(~input_layer[1917]),
      .e(~input_layer[1421]),
      .y(Y[1889]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1890_1
  function_67 neuron1890_1 (
      .a(input_layer[875]),
      .b(input_layer[2120]),
      .c(~input_layer[546]),
      .d(input_layer[1815]),
      .e(input_layer[1809]),
      .y(Y[1890]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1891_1
  function_104 neuron1891_1 (
      .a(input_layer[1607]),
      .b(~input_layer[1195]),
      .c(~input_layer[234]),
      .y(Y[1891]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_20 for neuron1892_1
  function_20 neuron1892_1 (
      .a(input_layer[1075]),
      .b(input_layer[1336]),
      .c(input_layer[955]),
      .d(~input_layer[1652]),
      .e(~input_layer[1357]),
      .f(input_layer[1226]),
      .y(Y[1892]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1893_1
  function_5 neuron1893_1 (
      .a(input_layer[1052]),
      .b(~input_layer[462]),
      .y(Y[1893]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1894_1
  function_188 neuron1894_1 (
      .a(input_layer[905]),
      .b(~input_layer[1499]),
      .c(~input_layer[1955]),
      .d(input_layer[417]),
      .e(input_layer[319]),
      .f(input_layer[2286]),
      .y(Y[1894]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1895_1
  function_10 neuron1895_1 (
      .a(input_layer[475]),
      .b(input_layer[113]),
      .c(~input_layer[1216]),
      .d(input_layer[1886]),
      .y(Y[1895]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_130 for neuron1896_1
  function_130 neuron1896_1 (
      .a(input_layer[682]),
      .b(input_layer[1703]),
      .c(input_layer[880]),
      .d(input_layer[358]),
      .e(~input_layer[36]),
      .f(input_layer[249]),
      .y(Y[1896]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_154 for neuron1897_1
  function_154 neuron1897_1 (
      .a(input_layer[552]),
      .b(input_layer[1791]),
      .c(~input_layer[2134]),
      .d(~input_layer[1967]),
      .e(input_layer[1421]),
      .y(Y[1897]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_139 for neuron1898_1
  function_139 neuron1898_1 (
      .a(input_layer[1553]),
      .b(~input_layer[519]),
      .c(input_layer[1679]),
      .d(~input_layer[1726]),
      .e(~input_layer[778]),
      .y(Y[1898]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1899_1
  function_16 neuron1899_1 (
      .a(~input_layer[351]),
      .b(input_layer[1844]),
      .c(input_layer[2206]),
      .y(Y[1899]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_166 for neuron1900_1
  function_166 neuron1900_1 (
      .a(~input_layer[1457]),
      .b(~input_layer[1604]),
      .c(input_layer[524]),
      .d(input_layer[1486]),
      .e(~input_layer[1180]),
      .f(input_layer[1261]),
      .y(Y[1900]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_421 for neuron1901_1
  function_421 neuron1901_1 (
      .a(~input_layer[1287]),
      .b(~input_layer[579]),
      .c(input_layer[641]),
      .d(~input_layer[1918]),
      .e(input_layer[1968]),
      .f(input_layer[1072]),
      .y(Y[1901]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1902_1
  function_107 neuron1902_1 (
      .a(~input_layer[1891]),
      .b(~input_layer[2063]),
      .c(input_layer[2126]),
      .d(~input_layer[319]),
      .y(Y[1902]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_143 for neuron1903_1
  function_143 neuron1903_1 (
      .a(input_layer[386]),
      .b(input_layer[455]),
      .c(input_layer[1667]),
      .d(~input_layer[1114]),
      .e(input_layer[1456]),
      .f(~input_layer[662]),
      .y(Y[1903]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1904_1
  function_11 neuron1904_1 (
      .a(input_layer[1567]),
      .b(input_layer[789]),
      .c(input_layer[1198]),
      .d(input_layer[1920]),
      .y(Y[1904]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_169 for neuron1905_1
  function_169 neuron1905_1 (
      .a(input_layer[1424]),
      .b(input_layer[1396]),
      .c(~input_layer[1297]),
      .d(~input_layer[1378]),
      .e(input_layer[662]),
      .f(~input_layer[1071]),
      .y(Y[1905]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_77 for neuron1906_1
  function_77 neuron1906_1 (
      .a(input_layer[2203]),
      .b(~input_layer[1947]),
      .c(input_layer[189]),
      .d(input_layer[1130]),
      .e(~input_layer[1495]),
      .f(input_layer[1275]),
      .y(Y[1906]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1907_1
  function_49 neuron1907_1 (
      .a(input_layer[1716]),
      .b(input_layer[461]),
      .c(~input_layer[1292]),
      .d(input_layer[112]),
      .e(input_layer[683]),
      .f(input_layer[2257]),
      .y(Y[1907]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_231 for neuron1908_1
  function_231 neuron1908_1 (
      .a(~input_layer[292]),
      .b(~input_layer[2226]),
      .c(~input_layer[2023]),
      .d(~input_layer[1473]),
      .e(input_layer[385]),
      .f(~input_layer[945]),
      .y(Y[1908]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1909_1
  function_16 neuron1909_1 (
      .a(input_layer[1475]),
      .b(input_layer[2081]),
      .c(input_layer[768]),
      .y(Y[1909]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_422 for neuron1910_1
  function_422 neuron1910_1 (
      .a(~input_layer[2074]),
      .b(input_layer[298]),
      .c(input_layer[217]),
      .d(~input_layer[1290]),
      .e(input_layer[267]),
      .f(~input_layer[1927]),
      .y(Y[1910]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1911_1
  function_11 neuron1911_1 (
      .a(input_layer[835]),
      .b(input_layer[482]),
      .c(input_layer[1013]),
      .d(~input_layer[1211]),
      .y(Y[1911]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_116 for neuron1912_1
  function_116 neuron1912_1 (
      .a(input_layer[2134]),
      .b(input_layer[1067]),
      .c(~input_layer[385]),
      .d(input_layer[2055]),
      .y(Y[1912]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_179 for neuron1913_1
  function_179 neuron1913_1 (
      .a(input_layer[657]),
      .b(~input_layer[1256]),
      .c(input_layer[882]),
      .d(input_layer[480]),
      .e(input_layer[2217]),
      .y(Y[1913]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_202 for neuron1914_1
  function_202 neuron1914_1 (
      .a(input_layer[1521]),
      .b(~input_layer[493]),
      .c(~input_layer[1633]),
      .d(input_layer[371]),
      .e(input_layer[611]),
      .y(Y[1914]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1915] = 1'b1;

  // instantiate function_142 for neuron1916_1
  function_142 neuron1916_1 (
      .a(~input_layer[2147]),
      .b(~input_layer[831]),
      .c(input_layer[292]),
      .d(input_layer[1189]),
      .e(input_layer[761]),
      .y(Y[1916]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_298 for neuron1917_1
  function_298 neuron1917_1 (
      .a(~input_layer[1194]),
      .b(input_layer[1725]),
      .c(input_layer[1413]),
      .d(~input_layer[1272]),
      .e(input_layer[2180]),
      .y(Y[1917]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_18 for neuron1918_1
  function_18 neuron1918_1 (
      .a(~input_layer[1823]),
      .b(~input_layer[551]),
      .c(~input_layer[320]),
      .d(~input_layer[413]),
      .e(input_layer[2063]),
      .y(Y[1918]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1919_1
  function_16 neuron1919_1 (
      .a(~input_layer[1962]),
      .b(input_layer[1524]),
      .c(input_layer[1079]),
      .y(Y[1919]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1920_1
  function_5 neuron1920_1 (
      .a(input_layer[229]),
      .b(input_layer[1650]),
      .y(Y[1920]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1921_1
  function_1 neuron1921_1 (
      .a(~input_layer[1454]),
      .b(~input_layer[1555]),
      .c(input_layer[1136]),
      .d(~input_layer[400]),
      .e(input_layer[463]),
      .f(~input_layer[529]),
      .y(Y[1921]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_67 for neuron1922_1
  function_67 neuron1922_1 (
      .a(input_layer[1585]),
      .b(input_layer[1072]),
      .c(~input_layer[531]),
      .d(input_layer[1744]),
      .e(~input_layer[299]),
      .y(Y[1922]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1923_1
  function_107 neuron1923_1 (
      .a(~input_layer[2311]),
      .b(~input_layer[1489]),
      .c(input_layer[869]),
      .d(~input_layer[1956]),
      .y(Y[1923]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1924_1
  function_25 neuron1924_1 (
      .a(input_layer[1918]),
      .b(input_layer[707]),
      .c(input_layer[2081]),
      .d(~input_layer[1050]),
      .e(input_layer[708]),
      .y(Y[1924]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_148 for neuron1925_1
  function_148 neuron1925_1 (
      .a(~input_layer[1993]),
      .b(input_layer[1292]),
      .c(input_layer[1287]),
      .d(~input_layer[596]),
      .y(Y[1925]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1926_1
  function_100 neuron1926_1 (
      .a(~input_layer[1464]),
      .b(input_layer[1572]),
      .c(input_layer[1620]),
      .y(Y[1926]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_423 for neuron1927_1
  function_423 neuron1927_1 (
      .a(~input_layer[488]),
      .b(input_layer[2217]),
      .c(input_layer[792]),
      .d(~input_layer[1703]),
      .e(input_layer[1981]),
      .f(~input_layer[1766]),
      .y(Y[1927]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_113 for neuron1928_1
  function_113 neuron1928_1 (
      .a(input_layer[1790]),
      .b(input_layer[763]),
      .c(input_layer[1686]),
      .d(input_layer[1734]),
      .e(input_layer[2335]),
      .f(~input_layer[643]),
      .y(Y[1928]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1929_1
  function_104 neuron1929_1 (
      .a(input_layer[1081]),
      .b(~input_layer[1215]),
      .c(~input_layer[2024]),
      .y(Y[1929]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1930_1
  function_54 neuron1930_1 (
      .a(input_layer[1998]),
      .b(input_layer[1507]),
      .c(input_layer[2330]),
      .d(~input_layer[555]),
      .e(input_layer[812]),
      .f(input_layer[374]),
      .y(Y[1930]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1931] = 1'b1;

  // instantiate function_125 for neuron1932_1
  function_125 neuron1932_1 (
      .a(~input_layer[550]),
      .b(~input_layer[374]),
      .c(input_layer[731]),
      .d(~input_layer[774]),
      .e(input_layer[1221]),
      .y(Y[1932]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1933_1
  function_3 neuron1933_1 (
      .a(input_layer[1070]),
      .b(input_layer[360]),
      .c(input_layer[2330]),
      .d(~input_layer[785]),
      .e(input_layer[468]),
      .y(Y[1933]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_93 for neuron1934_1
  function_93 neuron1934_1 (
      .a(~input_layer[1200]),
      .b(input_layer[1698]),
      .c(~input_layer[1749]),
      .d(~input_layer[2297]),
      .e(input_layer[1959]),
      .f(input_layer[2268]),
      .y(Y[1934]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_32 for neuron1935_1
  function_32 neuron1935_1 (
      .a(input_layer[1123]),
      .b(input_layer[1537]),
      .c(input_layer[1329]),
      .d(~input_layer[2201]),
      .y(Y[1935]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_3 for neuron1936_1
  function_3 neuron1936_1 (
      .a(input_layer[299]),
      .b(input_layer[218]),
      .c(~input_layer[1308]),
      .d(~input_layer[813]),
      .e(input_layer[2119]),
      .y(Y[1936]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1937_1
  function_12 neuron1937_1 (
      .a(~input_layer[2246]),
      .b(~input_layer[762]),
      .c(input_layer[981]),
      .y(Y[1937]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1938_1
  function_5 neuron1938_1 (
      .a(input_layer[1068]),
      .b(input_layer[1061]),
      .y(Y[1938]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1939_1
  function_1 neuron1939_1 (
      .a(~input_layer[751]),
      .b(~input_layer[1690]),
      .c(~input_layer[1270]),
      .d(~input_layer[1609]),
      .e(~input_layer[2095]),
      .f(~input_layer[2108]),
      .y(Y[1939]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_37 for neuron1940_1
  function_37 neuron1940_1 (
      .a(input_layer[743]),
      .b(input_layer[395]),
      .c(~input_layer[2217]),
      .d(~input_layer[1644]),
      .e(input_layer[1606]),
      .y(Y[1940]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1941_1
  function_12 neuron1941_1 (
      .a(~input_layer[1322]),
      .b(~input_layer[2324]),
      .c(~input_layer[1101]),
      .y(Y[1941]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1942_1
  function_35 neuron1942_1 (
      .a(~input_layer[1837]),
      .b(input_layer[2033]),
      .c(~input_layer[2307]),
      .d(~input_layer[1875]),
      .e(~input_layer[290]),
      .y(Y[1942]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1943_1
  function_11 neuron1943_1 (
      .a(input_layer[1625]),
      .b(input_layer[1371]),
      .c(input_layer[494]),
      .d(input_layer[559]),
      .y(Y[1943]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1944] = 1'b0;

  // instantiate function_67 for neuron1945_1
  function_67 neuron1945_1 (
      .a(input_layer[198]),
      .b(input_layer[2229]),
      .c(~input_layer[858]),
      .d(~input_layer[1170]),
      .e(input_layer[397]),
      .y(Y[1945]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_95 for neuron1946_1
  function_95 neuron1946_1 (
      .a(input_layer[1691]),
      .b(~input_layer[1335]),
      .c(input_layer[1325]),
      .d(~input_layer[1709]),
      .y(Y[1946]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_188 for neuron1947_1
  function_188 neuron1947_1 (
      .a(input_layer[1797]),
      .b(input_layer[826]),
      .c(input_layer[101]),
      .d(~input_layer[432]),
      .e(~input_layer[2012]),
      .f(~input_layer[1023]),
      .y(Y[1947]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_388 for neuron1948_1
  function_388 neuron1948_1 (
      .a(~input_layer[1707]),
      .b(~input_layer[1507]),
      .c(input_layer[1226]),
      .d(input_layer[1113]),
      .e(~input_layer[1748]),
      .y(Y[1948]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_5 for neuron1949_1
  function_5 neuron1949_1 (
      .a(input_layer[297]),
      .b(input_layer[462]),
      .y(Y[1949]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_107 for neuron1950_1
  function_107 neuron1950_1 (
      .a(~input_layer[1533]),
      .b(~input_layer[667]),
      .c(~input_layer[552]),
      .d(~input_layer[1947]),
      .y(Y[1950]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_21 for neuron1951_1
  function_21 neuron1951_1 (
      .a(~input_layer[2023]),
      .b(input_layer[471]),
      .c(~input_layer[1509]),
      .d(~input_layer[1406]),
      .y(Y[1951]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_1 for neuron1952_1
  function_1 neuron1952_1 (
      .a(~input_layer[825]),
      .b(~input_layer[1074]),
      .c(~input_layer[652]),
      .d(~input_layer[1539]),
      .e(~input_layer[1243]),
      .f(~input_layer[837]),
      .y(Y[1952]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1953_1
  function_11 neuron1953_1 (
      .a(input_layer[2071]),
      .b(input_layer[413]),
      .c(input_layer[1002]),
      .d(~input_layer[1555]),
      .y(Y[1953]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_192 for neuron1954_1
  function_192 neuron1954_1 (
      .a(~input_layer[1049]),
      .b(~input_layer[639]),
      .c(~input_layer[1133]),
      .d(input_layer[1060]),
      .e(~input_layer[523]),
      .f(~input_layer[489]),
      .y(Y[1954]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_35 for neuron1955_1
  function_35 neuron1955_1 (
      .a(~input_layer[1945]),
      .b(~input_layer[915]),
      .c(~input_layer[1928]),
      .d(input_layer[412]),
      .e(~input_layer[2177]),
      .y(Y[1955]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1956_1
  function_49 neuron1956_1 (
      .a(input_layer[984]),
      .b(input_layer[996]),
      .c(input_layer[456]),
      .d(~input_layer[392]),
      .e(input_layer[1422]),
      .f(input_layer[585]),
      .y(Y[1956]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_288 for neuron1957_1
  function_288 neuron1957_1 (
      .a(input_layer[2153]),
      .b(input_layer[222]),
      .c(~input_layer[2317]),
      .d(~input_layer[1696]),
      .e(input_layer[2142]),
      .f(~input_layer[838]),
      .y(Y[1957]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_125 for neuron1958_1
  function_125 neuron1958_1 (
      .a(~input_layer[277]),
      .b(input_layer[1286]),
      .c(~input_layer[2287]),
      .d(input_layer[1324]),
      .e(~input_layer[1233]),
      .y(Y[1958]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_196 for neuron1959_1
  function_196 neuron1959_1 (
      .a(input_layer[824]),
      .b(~input_layer[1471]),
      .c(input_layer[1971]),
      .d(~input_layer[925]),
      .e(input_layer[785]),
      .f(~input_layer[456]),
      .y(Y[1959]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_249 for neuron1960_1
  function_249 neuron1960_1 (
      .a(~input_layer[1421]),
      .b(input_layer[2029]),
      .c(input_layer[324]),
      .d(input_layer[678]),
      .e(~input_layer[535]),
      .f(~input_layer[1357]),
      .y(Y[1960]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_254 for neuron1961_1
  function_254 neuron1961_1 (
      .a(~input_layer[312]),
      .b(~input_layer[1168]),
      .c(~input_layer[1540]),
      .d(~input_layer[1498]),
      .e(input_layer[1818]),
      .f(input_layer[691]),
      .y(Y[1961]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_424 for neuron1962_1
  function_424 neuron1962_1 (
      .a(~input_layer[403]),
      .b(input_layer[1944]),
      .c(~input_layer[987]),
      .d(input_layer[1006]),
      .e(input_layer[145]),
      .f(input_layer[2053]),
      .y(Y[1962]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_224 for neuron1963_1
  function_224 neuron1963_1 (
      .a(input_layer[1019]),
      .b(~input_layer[287]),
      .c(~input_layer[1415]),
      .d(~input_layer[1042]),
      .y(Y[1963]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_306 for neuron1964_1
  function_306 neuron1964_1 (
      .a(input_layer[1744]),
      .b(~input_layer[1063]),
      .c(input_layer[1791]),
      .d(input_layer[1613]),
      .e(input_layer[2055]),
      .f(input_layer[670]),
      .y(Y[1964]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_33 for neuron1965_1
  function_33 neuron1965_1 (
      .a(~input_layer[1395]),
      .b(input_layer[1787]),
      .c(~input_layer[238]),
      .d(~input_layer[914]),
      .e(~input_layer[2197]),
      .y(Y[1965]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1966_1
  function_10 neuron1966_1 (
      .a(input_layer[317]),
      .b(input_layer[183]),
      .c(input_layer[529]),
      .d(~input_layer[2323]),
      .y(Y[1966]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_11 for neuron1967_1
  function_11 neuron1967_1 (
      .a(input_layer[485]),
      .b(input_layer[1414]),
      .c(input_layer[1419]),
      .d(~input_layer[879]),
      .y(Y[1967]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_117 for neuron1968_1
  function_117 neuron1968_1 (
      .a(~input_layer[2210]),
      .b(input_layer[1411]),
      .c(~input_layer[1752]),
      .d(~input_layer[1755]),
      .e(input_layer[1550]),
      .f(~input_layer[1011]),
      .y(Y[1968]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1969_1
  function_10 neuron1969_1 (
      .a(input_layer[1453]),
      .b(input_layer[599]),
      .c(~input_layer[1389]),
      .d(input_layer[779]),
      .y(Y[1969]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1970_1
  function_100 neuron1970_1 (
      .a(input_layer[130]),
      .b(~input_layer[1579]),
      .c(input_layer[1212]),
      .y(Y[1970]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1971_1
  function_12 neuron1971_1 (
      .a(~input_layer[1463]),
      .b(~input_layer[1558]),
      .c(input_layer[1237]),
      .y(Y[1971]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_425 for neuron1972_1
  function_425 neuron1972_1 (
      .a(~input_layer[1574]),
      .b(~input_layer[549]),
      .c(input_layer[1152]),
      .d(input_layer[1727]),
      .e(~input_layer[1944]),
      .f(input_layer[1279]),
      .y(Y[1972]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1973_1
  function_104 neuron1973_1 (
      .a(input_layer[2177]),
      .b(~input_layer[1480]),
      .c(~input_layer[908]),
      .y(Y[1973]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_10 for neuron1974_1
  function_10 neuron1974_1 (
      .a(input_layer[2224]),
      .b(input_layer[1778]),
      .c(~input_layer[1140]),
      .d(input_layer[2089]),
      .y(Y[1974]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_25 for neuron1975_1
  function_25 neuron1975_1 (
      .a(input_layer[1392]),
      .b(input_layer[1417]),
      .c(input_layer[112]),
      .d(input_layer[775]),
      .e(~input_layer[1822]),
      .y(Y[1975]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1976_1
  function_162 neuron1976_1 (
      .a(~input_layer[833]),
      .b(~input_layer[1011]),
      .c(input_layer[1651]),
      .d(~input_layer[1217]),
      .e(~input_layer[864]),
      .y(Y[1976]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_19 for neuron1977_1
  function_19 neuron1977_1 (
      .a(~input_layer[631]),
      .b(input_layer[2307]),
      .c(~input_layer[2134]),
      .d(~input_layer[1209]),
      .y(Y[1977]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_426 for neuron1978_1
  function_426 neuron1978_1 (
      .a(input_layer[718]),
      .b(input_layer[2242]),
      .c(~input_layer[1163]),
      .d(input_layer[1357]),
      .e(input_layer[1699]),
      .f(~input_layer[154]),
      .y(Y[1978]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1979_1
  function_64 neuron1979_1 (
      .a(~input_layer[1184]),
      .b(input_layer[320]),
      .c(input_layer[1494]),
      .d(input_layer[2258]),
      .e(~input_layer[1180]),
      .y(Y[1979]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_49 for neuron1980_1
  function_49 neuron1980_1 (
      .a(input_layer[608]),
      .b(input_layer[220]),
      .c(input_layer[752]),
      .d(input_layer[359]),
      .e(~input_layer[1115]),
      .f(input_layer[451]),
      .y(Y[1980]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_162 for neuron1981_1
  function_162 neuron1981_1 (
      .a(~input_layer[1400]),
      .b(~input_layer[2227]),
      .c(~input_layer[1185]),
      .d(input_layer[2075]),
      .e(~input_layer[2333]),
      .y(Y[1981]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_63 for neuron1982_1
  function_63 neuron1982_1 (
      .a(input_layer[556]),
      .b(input_layer[345]),
      .c(~input_layer[1356]),
      .d(input_layer[1816]),
      .y(Y[1982]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_404 for neuron1983_1
  function_404 neuron1983_1 (
      .a(~input_layer[1122]),
      .b(~input_layer[1529]),
      .c(input_layer[1300]),
      .d(~input_layer[289]),
      .e(input_layer[1083]),
      .f(~input_layer[603]),
      .y(Y[1983]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_115 for neuron1984_1
  function_115 neuron1984_1 (
      .a(input_layer[2206]),
      .b(~input_layer[781]),
      .c(~input_layer[2248]),
      .d(input_layer[133]),
      .e(input_layer[258]),
      .y(Y[1984]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_64 for neuron1985_1
  function_64 neuron1985_1 (
      .a(input_layer[1297]),
      .b(input_layer[279]),
      .c(input_layer[1954]),
      .d(input_layer[154]),
      .e(~input_layer[648]),
      .y(Y[1985]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_99 for neuron1986_1
  function_99 neuron1986_1 (
      .a(input_layer[1861]),
      .b(~input_layer[273]),
      .c(input_layer[1087]),
      .d(input_layer[1046]),
      .e(~input_layer[1206]),
      .f(~input_layer[2132]),
      .y(Y[1986]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_104 for neuron1987_1
  function_104 neuron1987_1 (
      .a(input_layer[2170]),
      .b(~input_layer[1558]),
      .c(~input_layer[1256]),
      .y(Y[1987]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_22 for neuron1988_1
  function_22 neuron1988_1 (
      .a(~input_layer[655]),
      .b(~input_layer[1950]),
      .c(~input_layer[1913]),
      .d(~input_layer[1994]),
      .e(input_layer[2198]),
      .f(~input_layer[1977]),
      .y(Y[1988]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_283 for neuron1989_1
  function_283 neuron1989_1 (
      .a(input_layer[1158]),
      .b(~input_layer[280]),
      .c(~input_layer[517]),
      .d(input_layer[2178]),
      .e(~input_layer[1678]),
      .f(~input_layer[337]),
      .y(Y[1989]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_100 for neuron1990_1
  function_100 neuron1990_1 (
      .a(input_layer[553]),
      .b(input_layer[1375]),
      .c(~input_layer[510]),
      .y(Y[1990]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_54 for neuron1991_1
  function_54 neuron1991_1 (
      .a(input_layer[977]),
      .b(input_layer[2216]),
      .c(~input_layer[1551]),
      .d(input_layer[328]),
      .e(input_layer[686]),
      .f(input_layer[545]),
      .y(Y[1991]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_45 for neuron1992_1
  function_45 neuron1992_1 (
      .a(~input_layer[228]),
      .b(input_layer[1220]),
      .c(~input_layer[1435]),
      .d(~input_layer[1256]),
      .e(~input_layer[400]),
      .f(~input_layer[1599]),
      .y(Y[1992]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_12 for neuron1993_1
  function_12 neuron1993_1 (
      .a(~input_layer[783]),
      .b(~input_layer[2042]),
      .c(~input_layer[877]),
      .y(Y[1993]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_348 for neuron1994_1
  function_348 neuron1994_1 (
      .a(~input_layer[1190]),
      .b(input_layer[683]),
      .c(input_layer[508]),
      .d(input_layer[155]),
      .e(~input_layer[840]),
      .f(~input_layer[208]),
      .y(Y[1994]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_204 for neuron1995_1
  function_204 neuron1995_1 (
      .a(~input_layer[930]),
      .b(input_layer[951]),
      .c(input_layer[2242]),
      .d(input_layer[596]),
      .e(input_layer[1138]),
      .y(Y[1995]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_61 for neuron1996_1
  function_61 neuron1996_1 (
      .a(~input_layer[365]),
      .b(~input_layer[1427]),
      .c(~input_layer[2065]),
      .d(input_layer[1831]),
      .e(input_layer[921]),
      .y(Y[1996]),
      .clk(clk),
      .rst(rst)
  );

  assign Y[1997] = 1'b1;

  // instantiate function_146 for neuron1998_1
  function_146 neuron1998_1 (
      .a(input_layer[1026]),
      .b(input_layer[2000]),
      .c(input_layer[668]),
      .d(~input_layer[2027]),
      .e(~input_layer[1195]),
      .y(Y[1998]),
      .clk(clk),
      .rst(rst)
  );

  // instantiate function_16 for neuron1999_1
  function_16 neuron1999_1 (
      .a(input_layer[1490]),
      .b(input_layer[417]),
      .c(input_layer[1579]),
      .y(Y[1999]),
      .clk(clk),
      .rst(rst)
  );

// total zero consts: 15
// total one  consts: 11
// total instantiations: 1974

  // Warning: Z[0] not driven (layer 3)
  // Warning: Z[1] not driven (layer 3)
  // Warning: Z[2] not driven (layer 3)
  // Warning: Z[3] not driven (layer 3)
  // Warning: Z[4] not driven (layer 3)
  // Warning: Z[5] not driven (layer 3)
  // Warning: Z[6] not driven (layer 3)
  // Warning: Z[7] not driven (layer 3)
  // Warning: Z[8] not driven (layer 3)
  // Warning: Z[9] not driven (layer 3)
  // Warning: Z[10] not driven (layer 3)
  // Warning: Z[11] not driven (layer 3)
  // Warning: Z[12] not driven (layer 3)
  // Warning: Z[13] not driven (layer 3)
  // Warning: Z[14] not driven (layer 3)
  // Warning: Z[15] not driven (layer 3)
  // Warning: Z[16] not driven (layer 3)
  // Warning: Z[17] not driven (layer 3)
  // Warning: Z[18] not driven (layer 3)
  // Warning: Z[19] not driven (layer 3)
  // Warning: Z[20] not driven (layer 3)
  // Warning: Z[21] not driven (layer 3)
  // Warning: Z[22] not driven (layer 3)
  // Warning: Z[23] not driven (layer 3)
  // Warning: Z[24] not driven (layer 3)
  // Warning: Z[25] not driven (layer 3)
  // Warning: Z[26] not driven (layer 3)
  // Warning: Z[27] not driven (layer 3)
  // Warning: Z[28] not driven (layer 3)
  // Warning: Z[29] not driven (layer 3)
  // Warning: Z[30] not driven (layer 3)
  // Warning: Z[31] not driven (layer 3)
  // Warning: Z[32] not driven (layer 3)
  // Warning: Z[33] not driven (layer 3)
  // Warning: Z[34] not driven (layer 3)
  // Warning: Z[35] not driven (layer 3)
  // Warning: Z[36] not driven (layer 3)
  // Warning: Z[37] not driven (layer 3)
  // Warning: Z[38] not driven (layer 3)
  // Warning: Z[39] not driven (layer 3)
  // Warning: Z[40] not driven (layer 3)
  // Warning: Z[41] not driven (layer 3)
  // Warning: Z[42] not driven (layer 3)
  // Warning: Z[43] not driven (layer 3)
  // Warning: Z[44] not driven (layer 3)
  // Warning: Z[45] not driven (layer 3)
  // Warning: Z[46] not driven (layer 3)
  // Warning: Z[47] not driven (layer 3)
  // Warning: Z[48] not driven (layer 3)
  // Warning: Z[49] not driven (layer 3)
  // Warning: Z[50] not driven (layer 3)
  // Warning: Z[51] not driven (layer 3)
  // Warning: Z[52] not driven (layer 3)
  // Warning: Z[53] not driven (layer 3)
  // Warning: Z[54] not driven (layer 3)
  // Warning: Z[55] not driven (layer 3)
  // Warning: Z[56] not driven (layer 3)
  // Warning: Z[57] not driven (layer 3)
  // Warning: Z[58] not driven (layer 3)
  // Warning: Z[59] not driven (layer 3)
  // Warning: Z[60] not driven (layer 3)
  // Warning: Z[61] not driven (layer 3)
  // Warning: Z[62] not driven (layer 3)
  // Warning: Z[63] not driven (layer 3)
  // Warning: Z[64] not driven (layer 3)
  // Warning: Z[65] not driven (layer 3)
  // Warning: Z[66] not driven (layer 3)
  // Warning: Z[67] not driven (layer 3)
  // Warning: Z[68] not driven (layer 3)
  // Warning: Z[69] not driven (layer 3)
  // Warning: Z[70] not driven (layer 3)
  // Warning: Z[71] not driven (layer 3)
  // Warning: Z[72] not driven (layer 3)
  // Warning: Z[73] not driven (layer 3)
  // Warning: Z[74] not driven (layer 3)
  // Warning: Z[75] not driven (layer 3)
  // Warning: Z[76] not driven (layer 3)
  // Warning: Z[77] not driven (layer 3)
  // Warning: Z[78] not driven (layer 3)
  // Warning: Z[79] not driven (layer 3)
  // Warning: Z[80] not driven (layer 3)
  // Warning: Z[81] not driven (layer 3)
  // Warning: Z[82] not driven (layer 3)
  // Warning: Z[83] not driven (layer 3)
  // Warning: Z[84] not driven (layer 3)
  // Warning: Z[85] not driven (layer 3)
  // Warning: Z[86] not driven (layer 3)
  // Warning: Z[87] not driven (layer 3)
  // Warning: Z[88] not driven (layer 3)
  // Warning: Z[89] not driven (layer 3)
  // Warning: Z[90] not driven (layer 3)
  // Warning: Z[91] not driven (layer 3)
  // Warning: Z[92] not driven (layer 3)
  // Warning: Z[93] not driven (layer 3)
  // Warning: Z[94] not driven (layer 3)
  // Warning: Z[95] not driven (layer 3)
  // Warning: Z[96] not driven (layer 3)
  // Warning: Z[97] not driven (layer 3)
  // Warning: Z[98] not driven (layer 3)
  // Warning: Z[99] not driven (layer 3)
  // Warning: Z[100] not driven (layer 3)
  // Warning: Z[101] not driven (layer 3)
  // Warning: Z[102] not driven (layer 3)
  // Warning: Z[103] not driven (layer 3)
  // Warning: Z[104] not driven (layer 3)
  // Warning: Z[105] not driven (layer 3)
  // Warning: Z[106] not driven (layer 3)
  // Warning: Z[107] not driven (layer 3)
  // Warning: Z[108] not driven (layer 3)
  // Warning: Z[109] not driven (layer 3)
  // Warning: Z[110] not driven (layer 3)
  // Warning: Z[111] not driven (layer 3)
  // Warning: Z[112] not driven (layer 3)
  // Warning: Z[113] not driven (layer 3)
  // Warning: Z[114] not driven (layer 3)
  // Warning: Z[115] not driven (layer 3)
  // Warning: Z[116] not driven (layer 3)
  // Warning: Z[117] not driven (layer 3)
  // Warning: Z[118] not driven (layer 3)
  // Warning: Z[119] not driven (layer 3)
  // Warning: Z[120] not driven (layer 3)
  // Warning: Z[121] not driven (layer 3)
  // Warning: Z[122] not driven (layer 3)
  // Warning: Z[123] not driven (layer 3)
  // Warning: Z[124] not driven (layer 3)
  // Warning: Z[125] not driven (layer 3)
  // Warning: Z[126] not driven (layer 3)
  // Warning: Z[127] not driven (layer 3)
  // Warning: Z[128] not driven (layer 3)
  // Warning: Z[129] not driven (layer 3)
  // Warning: Z[130] not driven (layer 3)
  // Warning: Z[131] not driven (layer 3)
  // Warning: Z[132] not driven (layer 3)
  // Warning: Z[133] not driven (layer 3)
  // Warning: Z[134] not driven (layer 3)
  // Warning: Z[135] not driven (layer 3)
  // Warning: Z[136] not driven (layer 3)
  // Warning: Z[137] not driven (layer 3)
  // Warning: Z[138] not driven (layer 3)
  // Warning: Z[139] not driven (layer 3)
  // Warning: Z[140] not driven (layer 3)
  // Warning: Z[141] not driven (layer 3)
  // Warning: Z[142] not driven (layer 3)
  // Warning: Z[143] not driven (layer 3)
  // Warning: Z[144] not driven (layer 3)
  // Warning: Z[145] not driven (layer 3)
  // Warning: Z[146] not driven (layer 3)
  // Warning: Z[147] not driven (layer 3)
  // Warning: Z[148] not driven (layer 3)
  // Warning: Z[149] not driven (layer 3)
  // Warning: Z[150] not driven (layer 3)
  // Warning: Z[151] not driven (layer 3)
  // Warning: Z[152] not driven (layer 3)
  // Warning: Z[153] not driven (layer 3)
  // Warning: Z[154] not driven (layer 3)
  // Warning: Z[155] not driven (layer 3)
  // Warning: Z[156] not driven (layer 3)
  // Warning: Z[157] not driven (layer 3)
  // Warning: Z[158] not driven (layer 3)
  // Warning: Z[159] not driven (layer 3)
  // Warning: Z[160] not driven (layer 3)
  // Warning: Z[161] not driven (layer 3)
  // Warning: Z[162] not driven (layer 3)
  // Warning: Z[163] not driven (layer 3)
  // Warning: Z[164] not driven (layer 3)
  // Warning: Z[165] not driven (layer 3)
  // Warning: Z[166] not driven (layer 3)
  // Warning: Z[167] not driven (layer 3)
  // Warning: Z[168] not driven (layer 3)
  // Warning: Z[169] not driven (layer 3)
  // Warning: Z[170] not driven (layer 3)
  // Warning: Z[171] not driven (layer 3)
  // Warning: Z[172] not driven (layer 3)
  // Warning: Z[173] not driven (layer 3)
  // Warning: Z[174] not driven (layer 3)
  // Warning: Z[175] not driven (layer 3)
  // Warning: Z[176] not driven (layer 3)
  // Warning: Z[177] not driven (layer 3)
  // Warning: Z[178] not driven (layer 3)
  // Warning: Z[179] not driven (layer 3)
  // Warning: Z[180] not driven (layer 3)
  // Warning: Z[181] not driven (layer 3)
  // Warning: Z[182] not driven (layer 3)
  // Warning: Z[183] not driven (layer 3)
  // Warning: Z[184] not driven (layer 3)
  // Warning: Z[185] not driven (layer 3)
  // Warning: Z[186] not driven (layer 3)
  // Warning: Z[187] not driven (layer 3)
  // Warning: Z[188] not driven (layer 3)
  // Warning: Z[189] not driven (layer 3)
  // Warning: Z[190] not driven (layer 3)
  // Warning: Z[191] not driven (layer 3)
  // Warning: Z[192] not driven (layer 3)
  // Warning: Z[193] not driven (layer 3)
  // Warning: Z[194] not driven (layer 3)
  // Warning: Z[195] not driven (layer 3)
  // Warning: Z[196] not driven (layer 3)
  // Warning: Z[197] not driven (layer 3)
  // Warning: Z[198] not driven (layer 3)
  // Warning: Z[199] not driven (layer 3)
  // Warning: Z[200] not driven (layer 3)
  // Warning: Z[201] not driven (layer 3)
  // Warning: Z[202] not driven (layer 3)
  // Warning: Z[203] not driven (layer 3)
  // Warning: Z[204] not driven (layer 3)
  // Warning: Z[205] not driven (layer 3)
  // Warning: Z[206] not driven (layer 3)
  // Warning: Z[207] not driven (layer 3)
  // Warning: Z[208] not driven (layer 3)
  // Warning: Z[209] not driven (layer 3)
  // Warning: Z[210] not driven (layer 3)
  // Warning: Z[211] not driven (layer 3)
  // Warning: Z[212] not driven (layer 3)
  // Warning: Z[213] not driven (layer 3)
  // Warning: Z[214] not driven (layer 3)
  // Warning: Z[215] not driven (layer 3)
  // Warning: Z[216] not driven (layer 3)
  // Warning: Z[217] not driven (layer 3)
  // Warning: Z[218] not driven (layer 3)
  // Warning: Z[219] not driven (layer 3)
  // Warning: Z[220] not driven (layer 3)
  // Warning: Z[221] not driven (layer 3)
  // Warning: Z[222] not driven (layer 3)
  // Warning: Z[223] not driven (layer 3)
  // Warning: Z[224] not driven (layer 3)
  // Warning: Z[225] not driven (layer 3)
  // Warning: Z[226] not driven (layer 3)
  // Warning: Z[227] not driven (layer 3)
  // Warning: Z[228] not driven (layer 3)
  // Warning: Z[229] not driven (layer 3)
  // Warning: Z[230] not driven (layer 3)
  // Warning: Z[231] not driven (layer 3)
  // Warning: Z[232] not driven (layer 3)
  // Warning: Z[233] not driven (layer 3)
  // Warning: Z[234] not driven (layer 3)
  // Warning: Z[235] not driven (layer 3)
  // Warning: Z[236] not driven (layer 3)
  // Warning: Z[237] not driven (layer 3)
  // Warning: Z[238] not driven (layer 3)
  // Warning: Z[239] not driven (layer 3)
  // Warning: Z[240] not driven (layer 3)
  // Warning: Z[241] not driven (layer 3)
  // Warning: Z[242] not driven (layer 3)
  // Warning: Z[243] not driven (layer 3)
  // Warning: Z[244] not driven (layer 3)
  // Warning: Z[245] not driven (layer 3)
  // Warning: Z[246] not driven (layer 3)
  // Warning: Z[247] not driven (layer 3)
  // Warning: Z[248] not driven (layer 3)
  // Warning: Z[249] not driven (layer 3)
  // Warning: Z[250] not driven (layer 3)
  // Warning: Z[251] not driven (layer 3)
  // Warning: Z[252] not driven (layer 3)
  // Warning: Z[253] not driven (layer 3)
  // Warning: Z[254] not driven (layer 3)
  // Warning: Z[255] not driven (layer 3)

endmodule
